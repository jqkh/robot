// DE0Qsys.v

// Generated using ACDS version 13.0sp1 232 at 2023.12.21.01:46:20

`timescale 1 ps / 1 ps
module DE0Qsys (
		input  wire        clk_50m_clk,       //     clk_50m.clk
		input  wire        reset_reset_n,     //       reset.reset_n
		input  wire        areset_export,     //      areset.export
		output wire        locked_export,     //      locked.export
		output wire        phasedone_export,  //   phasedone.export
		output wire [11:0] sdram_wires_addr,  // sdram_wires.addr
		output wire [1:0]  sdram_wires_ba,    //            .ba
		output wire        sdram_wires_cas_n, //            .cas_n
		output wire        sdram_wires_cke,   //            .cke
		output wire        sdram_wires_cs_n,  //            .cs_n
		inout  wire [15:0] sdram_wires_dq,    //            .dq
		output wire [1:0]  sdram_wires_dqm,   //            .dqm
		output wire        sdram_wires_ras_n, //            .ras_n
		output wire        sdram_wires_we_n,  //            .we_n
		input  wire        uart0_rxd,         //       uart0.rxd
		output wire        uart0_txd,         //            .txd
		output wire        dram_clk_clk,      //    dram_clk.clk
		output wire [9:0]  led_export,        //         led.export
		input  wire [3:0]  sw_export,         //          sw.export
		input  wire        button1_export,    //     button1.export
		input  wire        button2_export,    //     button2.export
		output wire [7:0]  hex0_export,       //        hex0.export
		output wire [7:0]  hex1_export,       //        hex1.export
		output wire [7:0]  hex2_export,       //        hex2.export
		output wire [7:0]  hex3_export        //        hex3.export
	);

	wire          syspll_c0_clk;                                                                                    // syspll:c0 -> [APB:clk, APB_m0_translator:clk, APB_m0_translator_avalon_universal_master_0_agent:clk, APB_s0_translator:clk, APB_s0_translator_avalon_universal_slave_0_agent:clk, APB_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, addr_router:clk, addr_router_001:clk, addr_router_002:clk, addr_router_003:clk, addr_router_004:clk, burst_adapter:clk, burst_adapter_001:clk, button1:clk, button1_s1_translator:clk, button1_s1_translator_avalon_universal_slave_0_agent:clk, button1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, button2:clk, button2_s1_translator:clk, button2_s1_translator_avalon_universal_slave_0_agent:clk, button2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, cmd_xbar_demux:clk, cmd_xbar_demux_001:clk, cmd_xbar_demux_002:clk, cmd_xbar_demux_003:clk, cmd_xbar_demux_004:clk, cmd_xbar_mux:clk, cmd_xbar_mux_001:clk, cmd_xbar_mux_002:clk, cmd_xbar_mux_003:clk, crosser:in_clk, crosser_001:out_clk, dma:clk, dma_control_port_slave_translator:clk, dma_control_port_slave_translator_avalon_universal_slave_0_agent:clk, dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, dma_read_master_translator:clk, dma_read_master_translator_avalon_universal_master_0_agent:clk, dma_write_master_translator:clk, dma_write_master_translator_avalon_universal_master_0_agent:clk, hex0:clk, hex0_s1_translator:clk, hex0_s1_translator_avalon_universal_slave_0_agent:clk, hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, hex1:clk, hex1_s1_translator:clk, hex1_s1_translator_avalon_universal_slave_0_agent:clk, hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, hex2:clk, hex2_s1_translator:clk, hex2_s1_translator_avalon_universal_slave_0_agent:clk, hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, hex3:clk, hex3_s1_translator:clk, hex3_s1_translator_avalon_universal_slave_0_agent:clk, hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, id_router:clk, id_router_001:clk, id_router_002:clk, id_router_003:clk, id_router_005:clk, id_router_006:clk, id_router_007:clk, id_router_008:clk, id_router_009:clk, id_router_010:clk, id_router_011:clk, id_router_012:clk, id_router_013:clk, id_router_014:clk, id_router_015:clk, irq_mapper:clk, jtag_uart:clk, jtag_uart_avalon_jtag_slave_translator:clk, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:clk, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, led:clk, led_s1_translator:clk, led_s1_translator_avalon_universal_slave_0_agent:clk, led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, limiter:clk, limiter_001:clk, nios2cpu:clk, nios2cpu_data_master_translator:clk, nios2cpu_data_master_translator_avalon_universal_master_0_agent:clk, nios2cpu_instruction_master_translator:clk, nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:clk, nios2cpu_jtag_debug_module_translator:clk, nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:clk, nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, rsp_xbar_demux:clk, rsp_xbar_demux_001:clk, rsp_xbar_demux_002:clk, rsp_xbar_demux_003:clk, rsp_xbar_demux_005:clk, rsp_xbar_demux_006:clk, rsp_xbar_demux_007:clk, rsp_xbar_demux_008:clk, rsp_xbar_demux_009:clk, rsp_xbar_demux_010:clk, rsp_xbar_demux_011:clk, rsp_xbar_demux_012:clk, rsp_xbar_demux_013:clk, rsp_xbar_demux_014:clk, rsp_xbar_demux_015:clk, rsp_xbar_mux:clk, rsp_xbar_mux_001:clk, rsp_xbar_mux_002:clk, rsp_xbar_mux_003:clk, rsp_xbar_mux_004:clk, rst_controller_001:clk, sdram_ctrl:clk, sdram_ctrl_s1_translator:clk, sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:clk, sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, sw:clk, sw_s1_translator:clk, sw_s1_translator_avalon_universal_slave_0_agent:clk, sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, timer:clk, timer_s1_translator:clk, timer_s1_translator_avalon_universal_slave_0_agent:clk, timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, uart0:clk, uart0_s1_translator:clk, uart0_s1_translator_avalon_universal_slave_0_agent:clk, uart0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, width_adapter:clk, width_adapter_001:clk]
	wire          nios2cpu_instruction_master_waitrequest;                                                          // nios2cpu_instruction_master_translator:av_waitrequest -> nios2cpu:i_waitrequest
	wire   [25:0] nios2cpu_instruction_master_address;                                                              // nios2cpu:i_address -> nios2cpu_instruction_master_translator:av_address
	wire          nios2cpu_instruction_master_read;                                                                 // nios2cpu:i_read -> nios2cpu_instruction_master_translator:av_read
	wire   [31:0] nios2cpu_instruction_master_readdata;                                                             // nios2cpu_instruction_master_translator:av_readdata -> nios2cpu:i_readdata
	wire    [7:0] dma_write_master_burstcount;                                                                      // dma:write_burstcount -> dma_write_master_translator:av_burstcount
	wire          dma_write_master_waitrequest;                                                                     // dma_write_master_translator:av_waitrequest -> dma:write_waitrequest
	wire   [31:0] dma_write_master_writedata;                                                                       // dma:write_writedata -> dma_write_master_translator:av_writedata
	wire   [25:0] dma_write_master_address;                                                                         // dma:write_address -> dma_write_master_translator:av_address
	wire          dma_write_master_chipselect;                                                                      // dma:write_chipselect -> dma_write_master_translator:av_chipselect
	wire          dma_write_master_write;                                                                           // dma:write_write_n -> dma_write_master_translator:av_write
	wire    [3:0] dma_write_master_byteenable;                                                                      // dma:write_byteenable -> dma_write_master_translator:av_byteenable
	wire          nios2cpu_data_master_waitrequest;                                                                 // nios2cpu_data_master_translator:av_waitrequest -> nios2cpu:d_waitrequest
	wire   [31:0] nios2cpu_data_master_writedata;                                                                   // nios2cpu:d_writedata -> nios2cpu_data_master_translator:av_writedata
	wire   [25:0] nios2cpu_data_master_address;                                                                     // nios2cpu:d_address -> nios2cpu_data_master_translator:av_address
	wire          nios2cpu_data_master_write;                                                                       // nios2cpu:d_write -> nios2cpu_data_master_translator:av_write
	wire          nios2cpu_data_master_read;                                                                        // nios2cpu:d_read -> nios2cpu_data_master_translator:av_read
	wire   [31:0] nios2cpu_data_master_readdata;                                                                    // nios2cpu_data_master_translator:av_readdata -> nios2cpu:d_readdata
	wire          nios2cpu_data_master_debugaccess;                                                                 // nios2cpu:jtag_debug_module_debugaccess_to_roms -> nios2cpu_data_master_translator:av_debugaccess
	wire    [3:0] nios2cpu_data_master_byteenable;                                                                  // nios2cpu:d_byteenable -> nios2cpu_data_master_translator:av_byteenable
	wire    [7:0] dma_read_master_burstcount;                                                                       // dma:read_burstcount -> dma_read_master_translator:av_burstcount
	wire          dma_read_master_waitrequest;                                                                      // dma_read_master_translator:av_waitrequest -> dma:read_waitrequest
	wire   [25:0] dma_read_master_address;                                                                          // dma:read_address -> dma_read_master_translator:av_address
	wire          dma_read_master_chipselect;                                                                       // dma:read_chipselect -> dma_read_master_translator:av_chipselect
	wire          dma_read_master_read;                                                                             // dma:read_read_n -> dma_read_master_translator:av_read
	wire   [31:0] dma_read_master_readdata;                                                                         // dma_read_master_translator:av_readdata -> dma:read_readdata
	wire          dma_read_master_readdatavalid;                                                                    // dma_read_master_translator:av_readdatavalid -> dma:read_readdatavalid
	wire          nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest;                            // nios2cpu:jtag_debug_module_waitrequest -> nios2cpu_jtag_debug_module_translator:av_waitrequest
	wire   [31:0] nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                              // nios2cpu_jtag_debug_module_translator:av_writedata -> nios2cpu:jtag_debug_module_writedata
	wire    [8:0] nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_address;                                // nios2cpu_jtag_debug_module_translator:av_address -> nios2cpu:jtag_debug_module_address
	wire          nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_write;                                  // nios2cpu_jtag_debug_module_translator:av_write -> nios2cpu:jtag_debug_module_write
	wire          nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_read;                                   // nios2cpu_jtag_debug_module_translator:av_read -> nios2cpu:jtag_debug_module_read
	wire   [31:0] nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                               // nios2cpu:jtag_debug_module_readdata -> nios2cpu_jtag_debug_module_translator:av_readdata
	wire          nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                            // nios2cpu_jtag_debug_module_translator:av_debugaccess -> nios2cpu:jtag_debug_module_debugaccess
	wire    [3:0] nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                             // nios2cpu_jtag_debug_module_translator:av_byteenable -> nios2cpu:jtag_debug_module_byteenable
	wire          sdram_ctrl_s1_translator_avalon_anti_slave_0_waitrequest;                                         // sdram_ctrl:za_waitrequest -> sdram_ctrl_s1_translator:av_waitrequest
	wire   [15:0] sdram_ctrl_s1_translator_avalon_anti_slave_0_writedata;                                           // sdram_ctrl_s1_translator:av_writedata -> sdram_ctrl:az_data
	wire   [21:0] sdram_ctrl_s1_translator_avalon_anti_slave_0_address;                                             // sdram_ctrl_s1_translator:av_address -> sdram_ctrl:az_addr
	wire          sdram_ctrl_s1_translator_avalon_anti_slave_0_chipselect;                                          // sdram_ctrl_s1_translator:av_chipselect -> sdram_ctrl:az_cs
	wire          sdram_ctrl_s1_translator_avalon_anti_slave_0_write;                                               // sdram_ctrl_s1_translator:av_write -> sdram_ctrl:az_wr_n
	wire          sdram_ctrl_s1_translator_avalon_anti_slave_0_read;                                                // sdram_ctrl_s1_translator:av_read -> sdram_ctrl:az_rd_n
	wire   [15:0] sdram_ctrl_s1_translator_avalon_anti_slave_0_readdata;                                            // sdram_ctrl:za_data -> sdram_ctrl_s1_translator:av_readdata
	wire          sdram_ctrl_s1_translator_avalon_anti_slave_0_readdatavalid;                                       // sdram_ctrl:za_valid -> sdram_ctrl_s1_translator:av_readdatavalid
	wire    [1:0] sdram_ctrl_s1_translator_avalon_anti_slave_0_byteenable;                                          // sdram_ctrl_s1_translator:av_byteenable -> sdram_ctrl:az_be_n
	wire   [25:0] dma_control_port_slave_translator_avalon_anti_slave_0_writedata;                                  // dma_control_port_slave_translator:av_writedata -> dma:dma_ctl_writedata
	wire    [2:0] dma_control_port_slave_translator_avalon_anti_slave_0_address;                                    // dma_control_port_slave_translator:av_address -> dma:dma_ctl_address
	wire          dma_control_port_slave_translator_avalon_anti_slave_0_chipselect;                                 // dma_control_port_slave_translator:av_chipselect -> dma:dma_ctl_chipselect
	wire          dma_control_port_slave_translator_avalon_anti_slave_0_write;                                      // dma_control_port_slave_translator:av_write -> dma:dma_ctl_write_n
	wire   [25:0] dma_control_port_slave_translator_avalon_anti_slave_0_readdata;                                   // dma:dma_ctl_readdata -> dma_control_port_slave_translator:av_readdata
	wire          apb_s0_translator_avalon_anti_slave_0_waitrequest;                                                // APB:s0_waitrequest -> APB_s0_translator:av_waitrequest
	wire    [0:0] apb_s0_translator_avalon_anti_slave_0_burstcount;                                                 // APB_s0_translator:av_burstcount -> APB:s0_burstcount
	wire   [31:0] apb_s0_translator_avalon_anti_slave_0_writedata;                                                  // APB_s0_translator:av_writedata -> APB:s0_writedata
	wire    [9:0] apb_s0_translator_avalon_anti_slave_0_address;                                                    // APB_s0_translator:av_address -> APB:s0_address
	wire          apb_s0_translator_avalon_anti_slave_0_write;                                                      // APB_s0_translator:av_write -> APB:s0_write
	wire          apb_s0_translator_avalon_anti_slave_0_read;                                                       // APB_s0_translator:av_read -> APB:s0_read
	wire   [31:0] apb_s0_translator_avalon_anti_slave_0_readdata;                                                   // APB:s0_readdata -> APB_s0_translator:av_readdata
	wire          apb_s0_translator_avalon_anti_slave_0_debugaccess;                                                // APB_s0_translator:av_debugaccess -> APB:s0_debugaccess
	wire          apb_s0_translator_avalon_anti_slave_0_readdatavalid;                                              // APB:s0_readdatavalid -> APB_s0_translator:av_readdatavalid
	wire    [3:0] apb_s0_translator_avalon_anti_slave_0_byteenable;                                                 // APB_s0_translator:av_byteenable -> APB:s0_byteenable
	wire   [31:0] syspll_pll_slave_translator_avalon_anti_slave_0_writedata;                                        // syspll_pll_slave_translator:av_writedata -> syspll:writedata
	wire    [1:0] syspll_pll_slave_translator_avalon_anti_slave_0_address;                                          // syspll_pll_slave_translator:av_address -> syspll:address
	wire          syspll_pll_slave_translator_avalon_anti_slave_0_write;                                            // syspll_pll_slave_translator:av_write -> syspll:write
	wire          syspll_pll_slave_translator_avalon_anti_slave_0_read;                                             // syspll_pll_slave_translator:av_read -> syspll:read
	wire   [31:0] syspll_pll_slave_translator_avalon_anti_slave_0_readdata;                                         // syspll:readdata -> syspll_pll_slave_translator:av_readdata
	wire    [0:0] apb_m0_burstcount;                                                                                // APB:m0_burstcount -> APB_m0_translator:av_burstcount
	wire          apb_m0_waitrequest;                                                                               // APB_m0_translator:av_waitrequest -> APB:m0_waitrequest
	wire    [9:0] apb_m0_address;                                                                                   // APB:m0_address -> APB_m0_translator:av_address
	wire   [31:0] apb_m0_writedata;                                                                                 // APB:m0_writedata -> APB_m0_translator:av_writedata
	wire          apb_m0_write;                                                                                     // APB:m0_write -> APB_m0_translator:av_write
	wire          apb_m0_read;                                                                                      // APB:m0_read -> APB_m0_translator:av_read
	wire   [31:0] apb_m0_readdata;                                                                                  // APB_m0_translator:av_readdata -> APB:m0_readdata
	wire          apb_m0_debugaccess;                                                                               // APB:m0_debugaccess -> APB_m0_translator:av_debugaccess
	wire    [3:0] apb_m0_byteenable;                                                                                // APB:m0_byteenable -> APB_m0_translator:av_byteenable
	wire          apb_m0_readdatavalid;                                                                             // APB_m0_translator:av_readdatavalid -> APB:m0_readdatavalid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                           // jtag_uart:av_waitrequest -> jtag_uart_avalon_jtag_slave_translator:av_waitrequest
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                             // jtag_uart_avalon_jtag_slave_translator:av_writedata -> jtag_uart:av_writedata
	wire    [0:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                               // jtag_uart_avalon_jtag_slave_translator:av_address -> jtag_uart:av_address
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                            // jtag_uart_avalon_jtag_slave_translator:av_chipselect -> jtag_uart:av_chipselect
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                 // jtag_uart_avalon_jtag_slave_translator:av_write -> jtag_uart:av_write_n
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                  // jtag_uart_avalon_jtag_slave_translator:av_read -> jtag_uart:av_read_n
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                              // jtag_uart:av_readdata -> jtag_uart_avalon_jtag_slave_translator:av_readdata
	wire   [15:0] timer_s1_translator_avalon_anti_slave_0_writedata;                                                // timer_s1_translator:av_writedata -> timer:writedata
	wire    [2:0] timer_s1_translator_avalon_anti_slave_0_address;                                                  // timer_s1_translator:av_address -> timer:address
	wire          timer_s1_translator_avalon_anti_slave_0_chipselect;                                               // timer_s1_translator:av_chipselect -> timer:chipselect
	wire          timer_s1_translator_avalon_anti_slave_0_write;                                                    // timer_s1_translator:av_write -> timer:write_n
	wire   [15:0] timer_s1_translator_avalon_anti_slave_0_readdata;                                                 // timer:readdata -> timer_s1_translator:av_readdata
	wire   [15:0] uart0_s1_translator_avalon_anti_slave_0_writedata;                                                // uart0_s1_translator:av_writedata -> uart0:writedata
	wire    [2:0] uart0_s1_translator_avalon_anti_slave_0_address;                                                  // uart0_s1_translator:av_address -> uart0:address
	wire          uart0_s1_translator_avalon_anti_slave_0_chipselect;                                               // uart0_s1_translator:av_chipselect -> uart0:chipselect
	wire          uart0_s1_translator_avalon_anti_slave_0_write;                                                    // uart0_s1_translator:av_write -> uart0:write_n
	wire          uart0_s1_translator_avalon_anti_slave_0_read;                                                     // uart0_s1_translator:av_read -> uart0:read_n
	wire   [15:0] uart0_s1_translator_avalon_anti_slave_0_readdata;                                                 // uart0:readdata -> uart0_s1_translator:av_readdata
	wire          uart0_s1_translator_avalon_anti_slave_0_begintransfer;                                            // uart0_s1_translator:av_begintransfer -> uart0:begintransfer
	wire    [1:0] sw_s1_translator_avalon_anti_slave_0_address;                                                     // sw_s1_translator:av_address -> sw:address
	wire   [31:0] sw_s1_translator_avalon_anti_slave_0_readdata;                                                    // sw:readdata -> sw_s1_translator:av_readdata
	wire   [31:0] led_s1_translator_avalon_anti_slave_0_writedata;                                                  // led_s1_translator:av_writedata -> led:writedata
	wire    [1:0] led_s1_translator_avalon_anti_slave_0_address;                                                    // led_s1_translator:av_address -> led:address
	wire          led_s1_translator_avalon_anti_slave_0_chipselect;                                                 // led_s1_translator:av_chipselect -> led:chipselect
	wire          led_s1_translator_avalon_anti_slave_0_write;                                                      // led_s1_translator:av_write -> led:write_n
	wire   [31:0] led_s1_translator_avalon_anti_slave_0_readdata;                                                   // led:readdata -> led_s1_translator:av_readdata
	wire   [31:0] button1_s1_translator_avalon_anti_slave_0_writedata;                                              // button1_s1_translator:av_writedata -> button1:writedata
	wire    [1:0] button1_s1_translator_avalon_anti_slave_0_address;                                                // button1_s1_translator:av_address -> button1:address
	wire          button1_s1_translator_avalon_anti_slave_0_chipselect;                                             // button1_s1_translator:av_chipselect -> button1:chipselect
	wire          button1_s1_translator_avalon_anti_slave_0_write;                                                  // button1_s1_translator:av_write -> button1:write_n
	wire   [31:0] button1_s1_translator_avalon_anti_slave_0_readdata;                                               // button1:readdata -> button1_s1_translator:av_readdata
	wire    [1:0] button2_s1_translator_avalon_anti_slave_0_address;                                                // button2_s1_translator:av_address -> button2:address
	wire   [31:0] button2_s1_translator_avalon_anti_slave_0_readdata;                                               // button2:readdata -> button2_s1_translator:av_readdata
	wire   [31:0] hex0_s1_translator_avalon_anti_slave_0_writedata;                                                 // hex0_s1_translator:av_writedata -> hex0:writedata
	wire    [1:0] hex0_s1_translator_avalon_anti_slave_0_address;                                                   // hex0_s1_translator:av_address -> hex0:address
	wire          hex0_s1_translator_avalon_anti_slave_0_chipselect;                                                // hex0_s1_translator:av_chipselect -> hex0:chipselect
	wire          hex0_s1_translator_avalon_anti_slave_0_write;                                                     // hex0_s1_translator:av_write -> hex0:write_n
	wire   [31:0] hex0_s1_translator_avalon_anti_slave_0_readdata;                                                  // hex0:readdata -> hex0_s1_translator:av_readdata
	wire   [31:0] hex1_s1_translator_avalon_anti_slave_0_writedata;                                                 // hex1_s1_translator:av_writedata -> hex1:writedata
	wire    [1:0] hex1_s1_translator_avalon_anti_slave_0_address;                                                   // hex1_s1_translator:av_address -> hex1:address
	wire          hex1_s1_translator_avalon_anti_slave_0_chipselect;                                                // hex1_s1_translator:av_chipselect -> hex1:chipselect
	wire          hex1_s1_translator_avalon_anti_slave_0_write;                                                     // hex1_s1_translator:av_write -> hex1:write_n
	wire   [31:0] hex1_s1_translator_avalon_anti_slave_0_readdata;                                                  // hex1:readdata -> hex1_s1_translator:av_readdata
	wire   [31:0] hex2_s1_translator_avalon_anti_slave_0_writedata;                                                 // hex2_s1_translator:av_writedata -> hex2:writedata
	wire    [1:0] hex2_s1_translator_avalon_anti_slave_0_address;                                                   // hex2_s1_translator:av_address -> hex2:address
	wire          hex2_s1_translator_avalon_anti_slave_0_chipselect;                                                // hex2_s1_translator:av_chipselect -> hex2:chipselect
	wire          hex2_s1_translator_avalon_anti_slave_0_write;                                                     // hex2_s1_translator:av_write -> hex2:write_n
	wire   [31:0] hex2_s1_translator_avalon_anti_slave_0_readdata;                                                  // hex2:readdata -> hex2_s1_translator:av_readdata
	wire   [31:0] hex3_s1_translator_avalon_anti_slave_0_writedata;                                                 // hex3_s1_translator:av_writedata -> hex3:writedata
	wire    [1:0] hex3_s1_translator_avalon_anti_slave_0_address;                                                   // hex3_s1_translator:av_address -> hex3:address
	wire          hex3_s1_translator_avalon_anti_slave_0_chipselect;                                                // hex3_s1_translator:av_chipselect -> hex3:chipselect
	wire          hex3_s1_translator_avalon_anti_slave_0_write;                                                     // hex3_s1_translator:av_write -> hex3:write_n
	wire   [31:0] hex3_s1_translator_avalon_anti_slave_0_readdata;                                                  // hex3:readdata -> hex3_s1_translator:av_readdata
	wire          nios2cpu_instruction_master_translator_avalon_universal_master_0_waitrequest;                     // nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2cpu_instruction_master_translator:uav_waitrequest
	wire    [2:0] nios2cpu_instruction_master_translator_avalon_universal_master_0_burstcount;                      // nios2cpu_instruction_master_translator:uav_burstcount -> nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] nios2cpu_instruction_master_translator_avalon_universal_master_0_writedata;                       // nios2cpu_instruction_master_translator:uav_writedata -> nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [25:0] nios2cpu_instruction_master_translator_avalon_universal_master_0_address;                         // nios2cpu_instruction_master_translator:uav_address -> nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire          nios2cpu_instruction_master_translator_avalon_universal_master_0_lock;                            // nios2cpu_instruction_master_translator:uav_lock -> nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire          nios2cpu_instruction_master_translator_avalon_universal_master_0_write;                           // nios2cpu_instruction_master_translator:uav_write -> nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire          nios2cpu_instruction_master_translator_avalon_universal_master_0_read;                            // nios2cpu_instruction_master_translator:uav_read -> nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] nios2cpu_instruction_master_translator_avalon_universal_master_0_readdata;                        // nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2cpu_instruction_master_translator:uav_readdata
	wire          nios2cpu_instruction_master_translator_avalon_universal_master_0_debugaccess;                     // nios2cpu_instruction_master_translator:uav_debugaccess -> nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] nios2cpu_instruction_master_translator_avalon_universal_master_0_byteenable;                      // nios2cpu_instruction_master_translator:uav_byteenable -> nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          nios2cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid;                   // nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2cpu_instruction_master_translator:uav_readdatavalid
	wire          dma_write_master_translator_avalon_universal_master_0_waitrequest;                                // dma_write_master_translator_avalon_universal_master_0_agent:av_waitrequest -> dma_write_master_translator:uav_waitrequest
	wire    [9:0] dma_write_master_translator_avalon_universal_master_0_burstcount;                                 // dma_write_master_translator:uav_burstcount -> dma_write_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] dma_write_master_translator_avalon_universal_master_0_writedata;                                  // dma_write_master_translator:uav_writedata -> dma_write_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [25:0] dma_write_master_translator_avalon_universal_master_0_address;                                    // dma_write_master_translator:uav_address -> dma_write_master_translator_avalon_universal_master_0_agent:av_address
	wire          dma_write_master_translator_avalon_universal_master_0_lock;                                       // dma_write_master_translator:uav_lock -> dma_write_master_translator_avalon_universal_master_0_agent:av_lock
	wire          dma_write_master_translator_avalon_universal_master_0_write;                                      // dma_write_master_translator:uav_write -> dma_write_master_translator_avalon_universal_master_0_agent:av_write
	wire          dma_write_master_translator_avalon_universal_master_0_read;                                       // dma_write_master_translator:uav_read -> dma_write_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] dma_write_master_translator_avalon_universal_master_0_readdata;                                   // dma_write_master_translator_avalon_universal_master_0_agent:av_readdata -> dma_write_master_translator:uav_readdata
	wire          dma_write_master_translator_avalon_universal_master_0_debugaccess;                                // dma_write_master_translator:uav_debugaccess -> dma_write_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] dma_write_master_translator_avalon_universal_master_0_byteenable;                                 // dma_write_master_translator:uav_byteenable -> dma_write_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          dma_write_master_translator_avalon_universal_master_0_readdatavalid;                              // dma_write_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> dma_write_master_translator:uav_readdatavalid
	wire          nios2cpu_data_master_translator_avalon_universal_master_0_waitrequest;                            // nios2cpu_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2cpu_data_master_translator:uav_waitrequest
	wire    [2:0] nios2cpu_data_master_translator_avalon_universal_master_0_burstcount;                             // nios2cpu_data_master_translator:uav_burstcount -> nios2cpu_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] nios2cpu_data_master_translator_avalon_universal_master_0_writedata;                              // nios2cpu_data_master_translator:uav_writedata -> nios2cpu_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [25:0] nios2cpu_data_master_translator_avalon_universal_master_0_address;                                // nios2cpu_data_master_translator:uav_address -> nios2cpu_data_master_translator_avalon_universal_master_0_agent:av_address
	wire          nios2cpu_data_master_translator_avalon_universal_master_0_lock;                                   // nios2cpu_data_master_translator:uav_lock -> nios2cpu_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire          nios2cpu_data_master_translator_avalon_universal_master_0_write;                                  // nios2cpu_data_master_translator:uav_write -> nios2cpu_data_master_translator_avalon_universal_master_0_agent:av_write
	wire          nios2cpu_data_master_translator_avalon_universal_master_0_read;                                   // nios2cpu_data_master_translator:uav_read -> nios2cpu_data_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] nios2cpu_data_master_translator_avalon_universal_master_0_readdata;                               // nios2cpu_data_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2cpu_data_master_translator:uav_readdata
	wire          nios2cpu_data_master_translator_avalon_universal_master_0_debugaccess;                            // nios2cpu_data_master_translator:uav_debugaccess -> nios2cpu_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] nios2cpu_data_master_translator_avalon_universal_master_0_byteenable;                             // nios2cpu_data_master_translator:uav_byteenable -> nios2cpu_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          nios2cpu_data_master_translator_avalon_universal_master_0_readdatavalid;                          // nios2cpu_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2cpu_data_master_translator:uav_readdatavalid
	wire          dma_read_master_translator_avalon_universal_master_0_waitrequest;                                 // dma_read_master_translator_avalon_universal_master_0_agent:av_waitrequest -> dma_read_master_translator:uav_waitrequest
	wire    [9:0] dma_read_master_translator_avalon_universal_master_0_burstcount;                                  // dma_read_master_translator:uav_burstcount -> dma_read_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] dma_read_master_translator_avalon_universal_master_0_writedata;                                   // dma_read_master_translator:uav_writedata -> dma_read_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [25:0] dma_read_master_translator_avalon_universal_master_0_address;                                     // dma_read_master_translator:uav_address -> dma_read_master_translator_avalon_universal_master_0_agent:av_address
	wire          dma_read_master_translator_avalon_universal_master_0_lock;                                        // dma_read_master_translator:uav_lock -> dma_read_master_translator_avalon_universal_master_0_agent:av_lock
	wire          dma_read_master_translator_avalon_universal_master_0_write;                                       // dma_read_master_translator:uav_write -> dma_read_master_translator_avalon_universal_master_0_agent:av_write
	wire          dma_read_master_translator_avalon_universal_master_0_read;                                        // dma_read_master_translator:uav_read -> dma_read_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] dma_read_master_translator_avalon_universal_master_0_readdata;                                    // dma_read_master_translator_avalon_universal_master_0_agent:av_readdata -> dma_read_master_translator:uav_readdata
	wire          dma_read_master_translator_avalon_universal_master_0_debugaccess;                                 // dma_read_master_translator:uav_debugaccess -> dma_read_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] dma_read_master_translator_avalon_universal_master_0_byteenable;                                  // dma_read_master_translator:uav_byteenable -> dma_read_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          dma_read_master_translator_avalon_universal_master_0_readdatavalid;                               // dma_read_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> dma_read_master_translator:uav_readdatavalid
	wire          nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // nios2cpu_jtag_debug_module_translator:uav_waitrequest -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;               // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> nios2cpu_jtag_debug_module_translator:uav_burstcount
	wire   [31:0] nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> nios2cpu_jtag_debug_module_translator:uav_writedata
	wire   [25:0] nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                  // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> nios2cpu_jtag_debug_module_translator:uav_address
	wire          nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                    // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> nios2cpu_jtag_debug_module_translator:uav_write
	wire          nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                     // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> nios2cpu_jtag_debug_module_translator:uav_lock
	wire          nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                     // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> nios2cpu_jtag_debug_module_translator:uav_read
	wire   [31:0] nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                 // nios2cpu_jtag_debug_module_translator:uav_readdata -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // nios2cpu_jtag_debug_module_translator:uav_readdatavalid -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> nios2cpu_jtag_debug_module_translator:uav_debugaccess
	wire    [3:0] nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;               // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> nios2cpu_jtag_debug_module_translator:uav_byteenable
	wire          nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;             // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [106:0] nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;              // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;             // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [106:0] nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // sdram_ctrl_s1_translator:uav_waitrequest -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [1:0] sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sdram_ctrl_s1_translator:uav_burstcount
	wire   [15:0] sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sdram_ctrl_s1_translator:uav_writedata
	wire   [25:0] sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:m0_address -> sdram_ctrl_s1_translator:uav_address
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:m0_write -> sdram_ctrl_s1_translator:uav_write
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sdram_ctrl_s1_translator:uav_lock
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:m0_read -> sdram_ctrl_s1_translator:uav_read
	wire   [15:0] sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // sdram_ctrl_s1_translator:uav_readdata -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // sdram_ctrl_s1_translator:uav_readdatavalid -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sdram_ctrl_s1_translator:uav_debugaccess
	wire    [1:0] sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sdram_ctrl_s1_translator:uav_byteenable
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [88:0] sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [88:0] sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [17:0] sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                     // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [17:0] sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                      // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                     // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                  // dma_control_port_slave_translator:uav_waitrequest -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                   // dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> dma_control_port_slave_translator:uav_burstcount
	wire   [31:0] dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                    // dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> dma_control_port_slave_translator:uav_writedata
	wire   [25:0] dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_address;                      // dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_address -> dma_control_port_slave_translator:uav_address
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_write;                        // dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_write -> dma_control_port_slave_translator:uav_write
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_lock;                         // dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_lock -> dma_control_port_slave_translator:uav_lock
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_read;                         // dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_read -> dma_control_port_slave_translator:uav_read
	wire   [31:0] dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                     // dma_control_port_slave_translator:uav_readdata -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                // dma_control_port_slave_translator:uav_readdatavalid -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                  // dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> dma_control_port_slave_translator:uav_debugaccess
	wire    [3:0] dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                   // dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> dma_control_port_slave_translator:uav_byteenable
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;           // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                 // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;         // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [106:0] dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                  // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                 // dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;        // dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;              // dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;      // dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [106:0] dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;               // dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;              // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;            // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] dma_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;             // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;            // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          apb_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // APB_s0_translator:uav_waitrequest -> APB_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] apb_s0_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // APB_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> APB_s0_translator:uav_burstcount
	wire   [31:0] apb_s0_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // APB_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> APB_s0_translator:uav_writedata
	wire   [25:0] apb_s0_translator_avalon_universal_slave_0_agent_m0_address;                                      // APB_s0_translator_avalon_universal_slave_0_agent:m0_address -> APB_s0_translator:uav_address
	wire          apb_s0_translator_avalon_universal_slave_0_agent_m0_write;                                        // APB_s0_translator_avalon_universal_slave_0_agent:m0_write -> APB_s0_translator:uav_write
	wire          apb_s0_translator_avalon_universal_slave_0_agent_m0_lock;                                         // APB_s0_translator_avalon_universal_slave_0_agent:m0_lock -> APB_s0_translator:uav_lock
	wire          apb_s0_translator_avalon_universal_slave_0_agent_m0_read;                                         // APB_s0_translator_avalon_universal_slave_0_agent:m0_read -> APB_s0_translator:uav_read
	wire   [31:0] apb_s0_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // APB_s0_translator:uav_readdata -> APB_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          apb_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // APB_s0_translator:uav_readdatavalid -> APB_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          apb_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // APB_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> APB_s0_translator:uav_debugaccess
	wire    [3:0] apb_s0_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // APB_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> APB_s0_translator:uav_byteenable
	wire          apb_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // APB_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> APB_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          apb_s0_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // APB_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> APB_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          apb_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // APB_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> APB_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [106:0] apb_s0_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // APB_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> APB_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          apb_s0_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // APB_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> APB_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          apb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // APB_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> APB_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          apb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // APB_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> APB_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          apb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // APB_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> APB_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [106:0] apb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // APB_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> APB_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          apb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // APB_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> APB_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          apb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // APB_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> APB_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] apb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // APB_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> APB_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          apb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // APB_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> APB_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // syspll_pll_slave_translator:uav_waitrequest -> syspll_pll_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // syspll_pll_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> syspll_pll_slave_translator:uav_burstcount
	wire   [31:0] syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                          // syspll_pll_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> syspll_pll_slave_translator:uav_writedata
	wire   [25:0] syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_address;                            // syspll_pll_slave_translator_avalon_universal_slave_0_agent:m0_address -> syspll_pll_slave_translator:uav_address
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_write;                              // syspll_pll_slave_translator_avalon_universal_slave_0_agent:m0_write -> syspll_pll_slave_translator:uav_write
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock;                               // syspll_pll_slave_translator_avalon_universal_slave_0_agent:m0_lock -> syspll_pll_slave_translator:uav_lock
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_read;                               // syspll_pll_slave_translator_avalon_universal_slave_0_agent:m0_read -> syspll_pll_slave_translator:uav_read
	wire   [31:0] syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                           // syspll_pll_slave_translator:uav_readdata -> syspll_pll_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // syspll_pll_slave_translator:uav_readdatavalid -> syspll_pll_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // syspll_pll_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> syspll_pll_slave_translator:uav_debugaccess
	wire    [3:0] syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // syspll_pll_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> syspll_pll_slave_translator:uav_byteenable
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // syspll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // syspll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // syspll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [106:0] syspll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                        // syspll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> syspll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> syspll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> syspll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> syspll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [106:0] syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> syspll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // syspll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // syspll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // syspll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> syspll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                  // syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> syspll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                   // syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> syspll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                  // syspll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          apb_m0_translator_avalon_universal_master_0_waitrequest;                                          // APB_m0_translator_avalon_universal_master_0_agent:av_waitrequest -> APB_m0_translator:uav_waitrequest
	wire    [2:0] apb_m0_translator_avalon_universal_master_0_burstcount;                                           // APB_m0_translator:uav_burstcount -> APB_m0_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] apb_m0_translator_avalon_universal_master_0_writedata;                                            // APB_m0_translator:uav_writedata -> APB_m0_translator_avalon_universal_master_0_agent:av_writedata
	wire    [9:0] apb_m0_translator_avalon_universal_master_0_address;                                              // APB_m0_translator:uav_address -> APB_m0_translator_avalon_universal_master_0_agent:av_address
	wire          apb_m0_translator_avalon_universal_master_0_lock;                                                 // APB_m0_translator:uav_lock -> APB_m0_translator_avalon_universal_master_0_agent:av_lock
	wire          apb_m0_translator_avalon_universal_master_0_write;                                                // APB_m0_translator:uav_write -> APB_m0_translator_avalon_universal_master_0_agent:av_write
	wire          apb_m0_translator_avalon_universal_master_0_read;                                                 // APB_m0_translator:uav_read -> APB_m0_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] apb_m0_translator_avalon_universal_master_0_readdata;                                             // APB_m0_translator_avalon_universal_master_0_agent:av_readdata -> APB_m0_translator:uav_readdata
	wire          apb_m0_translator_avalon_universal_master_0_debugaccess;                                          // APB_m0_translator:uav_debugaccess -> APB_m0_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] apb_m0_translator_avalon_universal_master_0_byteenable;                                           // APB_m0_translator:uav_byteenable -> APB_m0_translator_avalon_universal_master_0_agent:av_byteenable
	wire          apb_m0_translator_avalon_universal_master_0_readdatavalid;                                        // APB_m0_translator_avalon_universal_master_0_agent:av_readdatavalid -> APB_m0_translator:uav_readdatavalid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // jtag_uart_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_avalon_jtag_slave_translator:uav_burstcount
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_avalon_jtag_slave_translator:uav_writedata
	wire    [9:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_avalon_jtag_slave_translator:uav_address
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_avalon_jtag_slave_translator:uav_write
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_avalon_jtag_slave_translator:uav_lock
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_avalon_jtag_slave_translator:uav_read
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // jtag_uart_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // jtag_uart_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_avalon_jtag_slave_translator:uav_debugaccess
	wire    [3:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_avalon_jtag_slave_translator:uav_byteenable
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [83:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [83:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // timer_s1_translator:uav_waitrequest -> timer_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // timer_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_s1_translator:uav_burstcount
	wire   [31:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // timer_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_s1_translator:uav_writedata
	wire    [9:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // timer_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_s1_translator:uav_address
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // timer_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_s1_translator:uav_write
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // timer_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_s1_translator:uav_lock
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // timer_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_s1_translator:uav_read
	wire   [31:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // timer_s1_translator:uav_readdata -> timer_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // timer_s1_translator:uav_readdatavalid -> timer_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // timer_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_s1_translator:uav_debugaccess
	wire    [3:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // timer_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_s1_translator:uav_byteenable
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // timer_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // timer_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // timer_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [83:0] timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // timer_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [83:0] timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          uart0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // uart0_s1_translator:uav_waitrequest -> uart0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] uart0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // uart0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> uart0_s1_translator:uav_burstcount
	wire   [31:0] uart0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // uart0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> uart0_s1_translator:uav_writedata
	wire    [9:0] uart0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // uart0_s1_translator_avalon_universal_slave_0_agent:m0_address -> uart0_s1_translator:uav_address
	wire          uart0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // uart0_s1_translator_avalon_universal_slave_0_agent:m0_write -> uart0_s1_translator:uav_write
	wire          uart0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // uart0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> uart0_s1_translator:uav_lock
	wire          uart0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // uart0_s1_translator_avalon_universal_slave_0_agent:m0_read -> uart0_s1_translator:uav_read
	wire   [31:0] uart0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // uart0_s1_translator:uav_readdata -> uart0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          uart0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // uart0_s1_translator:uav_readdatavalid -> uart0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          uart0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // uart0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> uart0_s1_translator:uav_debugaccess
	wire    [3:0] uart0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // uart0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> uart0_s1_translator:uav_byteenable
	wire          uart0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // uart0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> uart0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          uart0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // uart0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> uart0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          uart0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // uart0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> uart0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [83:0] uart0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // uart0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> uart0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          uart0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // uart0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> uart0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          uart0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // uart0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> uart0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          uart0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // uart0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> uart0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          uart0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // uart0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> uart0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [83:0] uart0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // uart0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> uart0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          uart0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // uart0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> uart0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          uart0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // uart0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> uart0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] uart0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // uart0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> uart0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          uart0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // uart0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> uart0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sw_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                   // sw_s1_translator:uav_waitrequest -> sw_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sw_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                    // sw_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sw_s1_translator:uav_burstcount
	wire   [31:0] sw_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                     // sw_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sw_s1_translator:uav_writedata
	wire    [9:0] sw_s1_translator_avalon_universal_slave_0_agent_m0_address;                                       // sw_s1_translator_avalon_universal_slave_0_agent:m0_address -> sw_s1_translator:uav_address
	wire          sw_s1_translator_avalon_universal_slave_0_agent_m0_write;                                         // sw_s1_translator_avalon_universal_slave_0_agent:m0_write -> sw_s1_translator:uav_write
	wire          sw_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                          // sw_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sw_s1_translator:uav_lock
	wire          sw_s1_translator_avalon_universal_slave_0_agent_m0_read;                                          // sw_s1_translator_avalon_universal_slave_0_agent:m0_read -> sw_s1_translator:uav_read
	wire   [31:0] sw_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                      // sw_s1_translator:uav_readdata -> sw_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sw_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                 // sw_s1_translator:uav_readdatavalid -> sw_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sw_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                   // sw_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sw_s1_translator:uav_debugaccess
	wire    [3:0] sw_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                    // sw_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sw_s1_translator:uav_byteenable
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                            // sw_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                  // sw_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                          // sw_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [83:0] sw_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                   // sw_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                  // sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sw_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                         // sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sw_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                               // sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sw_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                       // sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sw_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [83:0] sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                // sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sw_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                               // sw_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                             // sw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                              // sw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                             // sw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          led_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // led_s1_translator:uav_waitrequest -> led_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] led_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // led_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> led_s1_translator:uav_burstcount
	wire   [31:0] led_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // led_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> led_s1_translator:uav_writedata
	wire    [9:0] led_s1_translator_avalon_universal_slave_0_agent_m0_address;                                      // led_s1_translator_avalon_universal_slave_0_agent:m0_address -> led_s1_translator:uav_address
	wire          led_s1_translator_avalon_universal_slave_0_agent_m0_write;                                        // led_s1_translator_avalon_universal_slave_0_agent:m0_write -> led_s1_translator:uav_write
	wire          led_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                         // led_s1_translator_avalon_universal_slave_0_agent:m0_lock -> led_s1_translator:uav_lock
	wire          led_s1_translator_avalon_universal_slave_0_agent_m0_read;                                         // led_s1_translator_avalon_universal_slave_0_agent:m0_read -> led_s1_translator:uav_read
	wire   [31:0] led_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // led_s1_translator:uav_readdata -> led_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          led_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // led_s1_translator:uav_readdatavalid -> led_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          led_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // led_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> led_s1_translator:uav_debugaccess
	wire    [3:0] led_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // led_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> led_s1_translator:uav_byteenable
	wire          led_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // led_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          led_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // led_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          led_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // led_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [83:0] led_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // led_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          led_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> led_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> led_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> led_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> led_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [83:0] led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> led_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // led_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          button1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // button1_s1_translator:uav_waitrequest -> button1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] button1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // button1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> button1_s1_translator:uav_burstcount
	wire   [31:0] button1_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                // button1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> button1_s1_translator:uav_writedata
	wire    [9:0] button1_s1_translator_avalon_universal_slave_0_agent_m0_address;                                  // button1_s1_translator_avalon_universal_slave_0_agent:m0_address -> button1_s1_translator:uav_address
	wire          button1_s1_translator_avalon_universal_slave_0_agent_m0_write;                                    // button1_s1_translator_avalon_universal_slave_0_agent:m0_write -> button1_s1_translator:uav_write
	wire          button1_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                     // button1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> button1_s1_translator:uav_lock
	wire          button1_s1_translator_avalon_universal_slave_0_agent_m0_read;                                     // button1_s1_translator_avalon_universal_slave_0_agent:m0_read -> button1_s1_translator:uav_read
	wire   [31:0] button1_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // button1_s1_translator:uav_readdata -> button1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          button1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // button1_s1_translator:uav_readdatavalid -> button1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          button1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // button1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> button1_s1_translator:uav_debugaccess
	wire    [3:0] button1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // button1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> button1_s1_translator:uav_byteenable
	wire          button1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // button1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> button1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          button1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // button1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> button1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          button1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // button1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> button1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [83:0] button1_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                              // button1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> button1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          button1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // button1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> button1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          button1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // button1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> button1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          button1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // button1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> button1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          button1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // button1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> button1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [83:0] button1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // button1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> button1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          button1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // button1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> button1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          button1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // button1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> button1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] button1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // button1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> button1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          button1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // button1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> button1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          button2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // button2_s1_translator:uav_waitrequest -> button2_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] button2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // button2_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> button2_s1_translator:uav_burstcount
	wire   [31:0] button2_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                // button2_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> button2_s1_translator:uav_writedata
	wire    [9:0] button2_s1_translator_avalon_universal_slave_0_agent_m0_address;                                  // button2_s1_translator_avalon_universal_slave_0_agent:m0_address -> button2_s1_translator:uav_address
	wire          button2_s1_translator_avalon_universal_slave_0_agent_m0_write;                                    // button2_s1_translator_avalon_universal_slave_0_agent:m0_write -> button2_s1_translator:uav_write
	wire          button2_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                     // button2_s1_translator_avalon_universal_slave_0_agent:m0_lock -> button2_s1_translator:uav_lock
	wire          button2_s1_translator_avalon_universal_slave_0_agent_m0_read;                                     // button2_s1_translator_avalon_universal_slave_0_agent:m0_read -> button2_s1_translator:uav_read
	wire   [31:0] button2_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // button2_s1_translator:uav_readdata -> button2_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          button2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // button2_s1_translator:uav_readdatavalid -> button2_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          button2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // button2_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> button2_s1_translator:uav_debugaccess
	wire    [3:0] button2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // button2_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> button2_s1_translator:uav_byteenable
	wire          button2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // button2_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> button2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          button2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // button2_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> button2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          button2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // button2_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> button2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [83:0] button2_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                              // button2_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> button2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          button2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // button2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> button2_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          button2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // button2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> button2_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          button2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // button2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> button2_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          button2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // button2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> button2_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [83:0] button2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // button2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> button2_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          button2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // button2_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> button2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          button2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // button2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> button2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] button2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // button2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> button2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          button2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // button2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> button2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          hex0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // hex0_s1_translator:uav_waitrequest -> hex0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] hex0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // hex0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> hex0_s1_translator:uav_burstcount
	wire   [31:0] hex0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // hex0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> hex0_s1_translator:uav_writedata
	wire    [9:0] hex0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                     // hex0_s1_translator_avalon_universal_slave_0_agent:m0_address -> hex0_s1_translator:uav_address
	wire          hex0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                       // hex0_s1_translator_avalon_universal_slave_0_agent:m0_write -> hex0_s1_translator:uav_write
	wire          hex0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                        // hex0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> hex0_s1_translator:uav_lock
	wire          hex0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                        // hex0_s1_translator_avalon_universal_slave_0_agent:m0_read -> hex0_s1_translator:uav_read
	wire   [31:0] hex0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // hex0_s1_translator:uav_readdata -> hex0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          hex0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // hex0_s1_translator:uav_readdatavalid -> hex0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          hex0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // hex0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> hex0_s1_translator:uav_debugaccess
	wire    [3:0] hex0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // hex0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> hex0_s1_translator:uav_byteenable
	wire          hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // hex0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // hex0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // hex0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [83:0] hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // hex0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> hex0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> hex0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> hex0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> hex0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [83:0] hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> hex0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // hex0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          hex0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // hex0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> hex0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] hex0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // hex0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> hex0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          hex0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // hex0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> hex0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          hex1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // hex1_s1_translator:uav_waitrequest -> hex1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] hex1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // hex1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> hex1_s1_translator:uav_burstcount
	wire   [31:0] hex1_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // hex1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> hex1_s1_translator:uav_writedata
	wire    [9:0] hex1_s1_translator_avalon_universal_slave_0_agent_m0_address;                                     // hex1_s1_translator_avalon_universal_slave_0_agent:m0_address -> hex1_s1_translator:uav_address
	wire          hex1_s1_translator_avalon_universal_slave_0_agent_m0_write;                                       // hex1_s1_translator_avalon_universal_slave_0_agent:m0_write -> hex1_s1_translator:uav_write
	wire          hex1_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                        // hex1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> hex1_s1_translator:uav_lock
	wire          hex1_s1_translator_avalon_universal_slave_0_agent_m0_read;                                        // hex1_s1_translator_avalon_universal_slave_0_agent:m0_read -> hex1_s1_translator:uav_read
	wire   [31:0] hex1_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // hex1_s1_translator:uav_readdata -> hex1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          hex1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // hex1_s1_translator:uav_readdatavalid -> hex1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          hex1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // hex1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> hex1_s1_translator:uav_debugaccess
	wire    [3:0] hex1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // hex1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> hex1_s1_translator:uav_byteenable
	wire          hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // hex1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // hex1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // hex1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [83:0] hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // hex1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> hex1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> hex1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> hex1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> hex1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [83:0] hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> hex1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // hex1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          hex1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // hex1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> hex1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] hex1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // hex1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> hex1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          hex1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // hex1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> hex1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          hex2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // hex2_s1_translator:uav_waitrequest -> hex2_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] hex2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // hex2_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> hex2_s1_translator:uav_burstcount
	wire   [31:0] hex2_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // hex2_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> hex2_s1_translator:uav_writedata
	wire    [9:0] hex2_s1_translator_avalon_universal_slave_0_agent_m0_address;                                     // hex2_s1_translator_avalon_universal_slave_0_agent:m0_address -> hex2_s1_translator:uav_address
	wire          hex2_s1_translator_avalon_universal_slave_0_agent_m0_write;                                       // hex2_s1_translator_avalon_universal_slave_0_agent:m0_write -> hex2_s1_translator:uav_write
	wire          hex2_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                        // hex2_s1_translator_avalon_universal_slave_0_agent:m0_lock -> hex2_s1_translator:uav_lock
	wire          hex2_s1_translator_avalon_universal_slave_0_agent_m0_read;                                        // hex2_s1_translator_avalon_universal_slave_0_agent:m0_read -> hex2_s1_translator:uav_read
	wire   [31:0] hex2_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // hex2_s1_translator:uav_readdata -> hex2_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          hex2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // hex2_s1_translator:uav_readdatavalid -> hex2_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          hex2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // hex2_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> hex2_s1_translator:uav_debugaccess
	wire    [3:0] hex2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // hex2_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> hex2_s1_translator:uav_byteenable
	wire          hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // hex2_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // hex2_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // hex2_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [83:0] hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // hex2_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> hex2_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> hex2_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> hex2_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> hex2_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [83:0] hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> hex2_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // hex2_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          hex2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // hex2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> hex2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] hex2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // hex2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> hex2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          hex2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // hex2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> hex2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          hex3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // hex3_s1_translator:uav_waitrequest -> hex3_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] hex3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // hex3_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> hex3_s1_translator:uav_burstcount
	wire   [31:0] hex3_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // hex3_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> hex3_s1_translator:uav_writedata
	wire    [9:0] hex3_s1_translator_avalon_universal_slave_0_agent_m0_address;                                     // hex3_s1_translator_avalon_universal_slave_0_agent:m0_address -> hex3_s1_translator:uav_address
	wire          hex3_s1_translator_avalon_universal_slave_0_agent_m0_write;                                       // hex3_s1_translator_avalon_universal_slave_0_agent:m0_write -> hex3_s1_translator:uav_write
	wire          hex3_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                        // hex3_s1_translator_avalon_universal_slave_0_agent:m0_lock -> hex3_s1_translator:uav_lock
	wire          hex3_s1_translator_avalon_universal_slave_0_agent_m0_read;                                        // hex3_s1_translator_avalon_universal_slave_0_agent:m0_read -> hex3_s1_translator:uav_read
	wire   [31:0] hex3_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // hex3_s1_translator:uav_readdata -> hex3_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          hex3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // hex3_s1_translator:uav_readdatavalid -> hex3_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          hex3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // hex3_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> hex3_s1_translator:uav_debugaccess
	wire    [3:0] hex3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // hex3_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> hex3_s1_translator:uav_byteenable
	wire          hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // hex3_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // hex3_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // hex3_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [83:0] hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // hex3_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> hex3_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> hex3_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> hex3_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> hex3_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [83:0] hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> hex3_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // hex3_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          hex3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // hex3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> hex3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] hex3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // hex3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> hex3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          hex3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // hex3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> hex3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          nios2cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;            // nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          nios2cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                  // nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          nios2cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;          // nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [105:0] nios2cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                   // nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          nios2cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                  // addr_router:sink_ready -> nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          dma_write_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                       // dma_write_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          dma_write_master_translator_avalon_universal_master_0_agent_cp_valid;                             // dma_write_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire          dma_write_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                     // dma_write_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [105:0] dma_write_master_translator_avalon_universal_master_0_agent_cp_data;                              // dma_write_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire          dma_write_master_translator_avalon_universal_master_0_agent_cp_ready;                             // addr_router_001:sink_ready -> dma_write_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          nios2cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                   // nios2cpu_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	wire          nios2cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid;                         // nios2cpu_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	wire          nios2cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                 // nios2cpu_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	wire  [105:0] nios2cpu_data_master_translator_avalon_universal_master_0_agent_cp_data;                          // nios2cpu_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	wire          nios2cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready;                         // addr_router_002:sink_ready -> nios2cpu_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          dma_read_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                        // dma_read_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_003:sink_endofpacket
	wire          dma_read_master_translator_avalon_universal_master_0_agent_cp_valid;                              // dma_read_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_003:sink_valid
	wire          dma_read_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                      // dma_read_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_003:sink_startofpacket
	wire  [105:0] dma_read_master_translator_avalon_universal_master_0_agent_cp_data;                               // dma_read_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_003:sink_data
	wire          dma_read_master_translator_avalon_universal_master_0_agent_cp_ready;                              // addr_router_003:sink_ready -> dma_read_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire          nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                    // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire          nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [105:0] nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                     // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire          nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router:sink_ready -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire   [87:0] sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_001:sink_ready -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                  // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_valid;                        // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [105:0] dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_data;                         // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_ready;                        // id_router_002:sink_ready -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          apb_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // APB_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire          apb_s0_translator_avalon_universal_slave_0_agent_rp_valid;                                        // APB_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire          apb_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // APB_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [105:0] apb_s0_translator_avalon_universal_slave_0_agent_rp_data;                                         // APB_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire          apb_s0_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_003:sink_ready -> APB_s0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // syspll_pll_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid;                              // syspll_pll_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // syspll_pll_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [105:0] syspll_pll_slave_translator_avalon_universal_slave_0_agent_rp_data;                               // syspll_pll_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready;                              // id_router_004:sink_ready -> syspll_pll_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          apb_m0_translator_avalon_universal_master_0_agent_cp_endofpacket;                                 // APB_m0_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_004:sink_endofpacket
	wire          apb_m0_translator_avalon_universal_master_0_agent_cp_valid;                                       // APB_m0_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_004:sink_valid
	wire          apb_m0_translator_avalon_universal_master_0_agent_cp_startofpacket;                               // APB_m0_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_004:sink_startofpacket
	wire   [82:0] apb_m0_translator_avalon_universal_master_0_agent_cp_data;                                        // APB_m0_translator_avalon_universal_master_0_agent:cp_data -> addr_router_004:sink_data
	wire          apb_m0_translator_avalon_universal_master_0_agent_cp_ready;                                       // addr_router_004:sink_ready -> APB_m0_translator_avalon_universal_master_0_agent:cp_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire   [82:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_005:sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // timer_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // timer_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // timer_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire   [82:0] timer_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // timer_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_006:sink_ready -> timer_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          uart0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // uart0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire          uart0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // uart0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire          uart0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // uart0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire   [82:0] uart0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // uart0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire          uart0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_007:sink_ready -> uart0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                   // sw_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                         // sw_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                 // sw_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire   [82:0] sw_s1_translator_avalon_universal_slave_0_agent_rp_data;                                          // sw_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                         // id_router_008:sink_ready -> sw_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          led_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // led_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire          led_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                        // led_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire          led_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // led_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire   [82:0] led_s1_translator_avalon_universal_slave_0_agent_rp_data;                                         // led_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire          led_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_009:sink_ready -> led_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          button1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // button1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire          button1_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                    // button1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire          button1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // button1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire   [82:0] button1_s1_translator_avalon_universal_slave_0_agent_rp_data;                                     // button1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire          button1_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_010:sink_ready -> button1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          button2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // button2_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	wire          button2_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                    // button2_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	wire          button2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // button2_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	wire   [82:0] button2_s1_translator_avalon_universal_slave_0_agent_rp_data;                                     // button2_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	wire          button2_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_011:sink_ready -> button2_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          hex0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // hex0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	wire          hex0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                       // hex0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	wire          hex0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // hex0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	wire   [82:0] hex0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                        // hex0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	wire          hex0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_012:sink_ready -> hex0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          hex1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // hex1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	wire          hex1_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                       // hex1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	wire          hex1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // hex1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	wire   [82:0] hex1_s1_translator_avalon_universal_slave_0_agent_rp_data;                                        // hex1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	wire          hex1_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_013:sink_ready -> hex1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          hex2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // hex2_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_014:sink_endofpacket
	wire          hex2_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                       // hex2_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_014:sink_valid
	wire          hex2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // hex2_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_014:sink_startofpacket
	wire   [82:0] hex2_s1_translator_avalon_universal_slave_0_agent_rp_data;                                        // hex2_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_014:sink_data
	wire          hex2_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_014:sink_ready -> hex2_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          hex3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // hex3_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_015:sink_endofpacket
	wire          hex3_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                       // hex3_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_015:sink_valid
	wire          hex3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // hex3_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_015:sink_startofpacket
	wire   [82:0] hex3_s1_translator_avalon_universal_slave_0_agent_rp_data;                                        // hex3_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_015:sink_data
	wire          hex3_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_015:sink_ready -> hex3_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          addr_router_003_src_endofpacket;                                                                  // addr_router_003:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire          addr_router_003_src_valid;                                                                        // addr_router_003:src_valid -> limiter:cmd_sink_valid
	wire          addr_router_003_src_startofpacket;                                                                // addr_router_003:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [105:0] addr_router_003_src_data;                                                                         // addr_router_003:src_data -> limiter:cmd_sink_data
	wire    [4:0] addr_router_003_src_channel;                                                                      // addr_router_003:src_channel -> limiter:cmd_sink_channel
	wire          addr_router_003_src_ready;                                                                        // limiter:cmd_sink_ready -> addr_router_003:src_ready
	wire          limiter_rsp_src_endofpacket;                                                                      // limiter:rsp_src_endofpacket -> dma_read_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_rsp_src_valid;                                                                            // limiter:rsp_src_valid -> dma_read_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_rsp_src_startofpacket;                                                                    // limiter:rsp_src_startofpacket -> dma_read_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [105:0] limiter_rsp_src_data;                                                                             // limiter:rsp_src_data -> dma_read_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [4:0] limiter_rsp_src_channel;                                                                          // limiter:rsp_src_channel -> dma_read_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_rsp_src_ready;                                                                            // dma_read_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire          addr_router_004_src_endofpacket;                                                                  // addr_router_004:src_endofpacket -> limiter_001:cmd_sink_endofpacket
	wire          addr_router_004_src_valid;                                                                        // addr_router_004:src_valid -> limiter_001:cmd_sink_valid
	wire          addr_router_004_src_startofpacket;                                                                // addr_router_004:src_startofpacket -> limiter_001:cmd_sink_startofpacket
	wire   [82:0] addr_router_004_src_data;                                                                         // addr_router_004:src_data -> limiter_001:cmd_sink_data
	wire   [10:0] addr_router_004_src_channel;                                                                      // addr_router_004:src_channel -> limiter_001:cmd_sink_channel
	wire          addr_router_004_src_ready;                                                                        // limiter_001:cmd_sink_ready -> addr_router_004:src_ready
	wire          limiter_001_rsp_src_endofpacket;                                                                  // limiter_001:rsp_src_endofpacket -> APB_m0_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_001_rsp_src_valid;                                                                        // limiter_001:rsp_src_valid -> APB_m0_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_001_rsp_src_startofpacket;                                                                // limiter_001:rsp_src_startofpacket -> APB_m0_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [82:0] limiter_001_rsp_src_data;                                                                         // limiter_001:rsp_src_data -> APB_m0_translator_avalon_universal_master_0_agent:rp_data
	wire   [10:0] limiter_001_rsp_src_channel;                                                                      // limiter_001:rsp_src_channel -> APB_m0_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_001_rsp_src_ready;                                                                        // APB_m0_translator_avalon_universal_master_0_agent:rp_ready -> limiter_001:rsp_src_ready
	wire          burst_adapter_source0_endofpacket;                                                                // burst_adapter:source0_endofpacket -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_source0_valid;                                                                      // burst_adapter:source0_valid -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_source0_startofpacket;                                                              // burst_adapter:source0_startofpacket -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [87:0] burst_adapter_source0_data;                                                                       // burst_adapter:source0_data -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_source0_ready;                                                                      // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire    [4:0] burst_adapter_source0_channel;                                                                    // burst_adapter:source0_channel -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_001_source0_endofpacket;                                                            // burst_adapter_001:source0_endofpacket -> APB_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_001_source0_valid;                                                                  // burst_adapter_001:source0_valid -> APB_s0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_001_source0_startofpacket;                                                          // burst_adapter_001:source0_startofpacket -> APB_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [105:0] burst_adapter_001_source0_data;                                                                   // burst_adapter_001:source0_data -> APB_s0_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_001_source0_ready;                                                                  // APB_s0_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_001:source0_ready
	wire    [4:0] burst_adapter_001_source0_channel;                                                                // burst_adapter_001:source0_channel -> APB_s0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rst_controller_reset_out_reset;                                                                   // rst_controller:reset_out -> [crosser:out_reset, crosser_001:in_reset, id_router_004:reset, rsp_xbar_demux_004:reset, syspll:reset, syspll_pll_slave_translator:reset, syspll_pll_slave_translator_avalon_universal_slave_0_agent:reset, syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire          rst_controller_001_reset_out_reset;                                                               // rst_controller_001:reset_out -> [APB:reset, APB_m0_translator:reset, APB_m0_translator_avalon_universal_master_0_agent:reset, APB_s0_translator:reset, APB_s0_translator_avalon_universal_slave_0_agent:reset, APB_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router:reset, addr_router_001:reset, addr_router_002:reset, addr_router_003:reset, addr_router_004:reset, burst_adapter:reset, burst_adapter_001:reset, button1:reset_n, button1_s1_translator:reset, button1_s1_translator_avalon_universal_slave_0_agent:reset, button1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, button2:reset_n, button2_s1_translator:reset, button2_s1_translator_avalon_universal_slave_0_agent:reset, button2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_demux_002:reset, cmd_xbar_demux_003:reset, cmd_xbar_demux_004:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_002:reset, cmd_xbar_mux_003:reset, crosser:in_reset, crosser_001:out_reset, dma:system_reset_n, dma_control_port_slave_translator:reset, dma_control_port_slave_translator_avalon_universal_slave_0_agent:reset, dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, dma_read_master_translator:reset, dma_read_master_translator_avalon_universal_master_0_agent:reset, dma_write_master_translator:reset, dma_write_master_translator_avalon_universal_master_0_agent:reset, hex0:reset_n, hex0_s1_translator:reset, hex0_s1_translator_avalon_universal_slave_0_agent:reset, hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, hex1:reset_n, hex1_s1_translator:reset, hex1_s1_translator_avalon_universal_slave_0_agent:reset, hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, hex2:reset_n, hex2_s1_translator:reset, hex2_s1_translator_avalon_universal_slave_0_agent:reset, hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, hex3:reset_n, hex3_s1_translator:reset, hex3_s1_translator_avalon_universal_slave_0_agent:reset, hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, id_router_011:reset, id_router_012:reset, id_router_013:reset, id_router_014:reset, id_router_015:reset, irq_mapper:reset, jtag_uart:rst_n, jtag_uart_avalon_jtag_slave_translator:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, led:reset_n, led_s1_translator:reset, led_s1_translator_avalon_universal_slave_0_agent:reset, led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter:reset, limiter_001:reset, nios2cpu:reset_n, nios2cpu_data_master_translator:reset, nios2cpu_data_master_translator_avalon_universal_master_0_agent:reset, nios2cpu_instruction_master_translator:reset, nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:reset, nios2cpu_jtag_debug_module_translator:reset, nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_013:reset, rsp_xbar_demux_014:reset, rsp_xbar_demux_015:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, rsp_xbar_mux_002:reset, rsp_xbar_mux_003:reset, rsp_xbar_mux_004:reset, sdram_ctrl:reset_n, sdram_ctrl_s1_translator:reset, sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:reset, sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sw:reset_n, sw_s1_translator:reset, sw_s1_translator_avalon_universal_slave_0_agent:reset, sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer:reset_n, timer_s1_translator:reset, timer_s1_translator_avalon_universal_slave_0_agent:reset, timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, uart0:reset_n, uart0_s1_translator:reset, uart0_s1_translator_avalon_universal_slave_0_agent:reset, uart0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, width_adapter:reset, width_adapter_001:reset]
	wire          nios2cpu_jtag_debug_module_reset_reset;                                                           // nios2cpu:jtag_debug_module_resetrequest -> rst_controller_001:reset_in1
	wire          cmd_xbar_demux_src0_endofpacket;                                                                  // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                        // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                                // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [105:0] cmd_xbar_demux_src0_data;                                                                         // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire    [4:0] cmd_xbar_demux_src0_channel;                                                                      // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire          cmd_xbar_demux_src0_ready;                                                                        // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire          cmd_xbar_demux_src1_endofpacket;                                                                  // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire          cmd_xbar_demux_src1_valid;                                                                        // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire          cmd_xbar_demux_src1_startofpacket;                                                                // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [105:0] cmd_xbar_demux_src1_data;                                                                         // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire    [4:0] cmd_xbar_demux_src1_channel;                                                                      // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire          cmd_xbar_demux_src1_ready;                                                                        // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire          cmd_xbar_demux_src2_endofpacket;                                                                  // cmd_xbar_demux:src2_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	wire          cmd_xbar_demux_src2_valid;                                                                        // cmd_xbar_demux:src2_valid -> cmd_xbar_mux_002:sink0_valid
	wire          cmd_xbar_demux_src2_startofpacket;                                                                // cmd_xbar_demux:src2_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	wire  [105:0] cmd_xbar_demux_src2_data;                                                                         // cmd_xbar_demux:src2_data -> cmd_xbar_mux_002:sink0_data
	wire    [4:0] cmd_xbar_demux_src2_channel;                                                                      // cmd_xbar_demux:src2_channel -> cmd_xbar_mux_002:sink0_channel
	wire          cmd_xbar_demux_src2_ready;                                                                        // cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux:src2_ready
	wire          cmd_xbar_demux_src3_endofpacket;                                                                  // cmd_xbar_demux:src3_endofpacket -> cmd_xbar_mux_003:sink0_endofpacket
	wire          cmd_xbar_demux_src3_valid;                                                                        // cmd_xbar_demux:src3_valid -> cmd_xbar_mux_003:sink0_valid
	wire          cmd_xbar_demux_src3_startofpacket;                                                                // cmd_xbar_demux:src3_startofpacket -> cmd_xbar_mux_003:sink0_startofpacket
	wire  [105:0] cmd_xbar_demux_src3_data;                                                                         // cmd_xbar_demux:src3_data -> cmd_xbar_mux_003:sink0_data
	wire    [4:0] cmd_xbar_demux_src3_channel;                                                                      // cmd_xbar_demux:src3_channel -> cmd_xbar_mux_003:sink0_channel
	wire          cmd_xbar_demux_src3_ready;                                                                        // cmd_xbar_mux_003:sink0_ready -> cmd_xbar_demux:src3_ready
	wire          cmd_xbar_demux_001_src0_endofpacket;                                                              // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                                                    // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux_001:sink1_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                                            // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [105:0] cmd_xbar_demux_001_src0_data;                                                                     // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux_001:sink1_data
	wire    [4:0] cmd_xbar_demux_001_src0_channel;                                                                  // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux_001:sink1_channel
	wire          cmd_xbar_demux_001_src0_ready;                                                                    // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire          cmd_xbar_demux_001_src1_endofpacket;                                                              // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_003:sink1_endofpacket
	wire          cmd_xbar_demux_001_src1_valid;                                                                    // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_003:sink1_valid
	wire          cmd_xbar_demux_001_src1_startofpacket;                                                            // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_003:sink1_startofpacket
	wire  [105:0] cmd_xbar_demux_001_src1_data;                                                                     // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_003:sink1_data
	wire    [4:0] cmd_xbar_demux_001_src1_channel;                                                                  // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_003:sink1_channel
	wire          cmd_xbar_demux_001_src1_ready;                                                                    // cmd_xbar_mux_003:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire          cmd_xbar_demux_002_src0_endofpacket;                                                              // cmd_xbar_demux_002:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire          cmd_xbar_demux_002_src0_valid;                                                                    // cmd_xbar_demux_002:src0_valid -> cmd_xbar_mux:sink1_valid
	wire          cmd_xbar_demux_002_src0_startofpacket;                                                            // cmd_xbar_demux_002:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [105:0] cmd_xbar_demux_002_src0_data;                                                                     // cmd_xbar_demux_002:src0_data -> cmd_xbar_mux:sink1_data
	wire    [4:0] cmd_xbar_demux_002_src0_channel;                                                                  // cmd_xbar_demux_002:src0_channel -> cmd_xbar_mux:sink1_channel
	wire          cmd_xbar_demux_002_src0_ready;                                                                    // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_002:src0_ready
	wire          cmd_xbar_demux_002_src1_endofpacket;                                                              // cmd_xbar_demux_002:src1_endofpacket -> cmd_xbar_mux_001:sink2_endofpacket
	wire          cmd_xbar_demux_002_src1_valid;                                                                    // cmd_xbar_demux_002:src1_valid -> cmd_xbar_mux_001:sink2_valid
	wire          cmd_xbar_demux_002_src1_startofpacket;                                                            // cmd_xbar_demux_002:src1_startofpacket -> cmd_xbar_mux_001:sink2_startofpacket
	wire  [105:0] cmd_xbar_demux_002_src1_data;                                                                     // cmd_xbar_demux_002:src1_data -> cmd_xbar_mux_001:sink2_data
	wire    [4:0] cmd_xbar_demux_002_src1_channel;                                                                  // cmd_xbar_demux_002:src1_channel -> cmd_xbar_mux_001:sink2_channel
	wire          cmd_xbar_demux_002_src1_ready;                                                                    // cmd_xbar_mux_001:sink2_ready -> cmd_xbar_demux_002:src1_ready
	wire          cmd_xbar_demux_002_src2_endofpacket;                                                              // cmd_xbar_demux_002:src2_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	wire          cmd_xbar_demux_002_src2_valid;                                                                    // cmd_xbar_demux_002:src2_valid -> cmd_xbar_mux_002:sink1_valid
	wire          cmd_xbar_demux_002_src2_startofpacket;                                                            // cmd_xbar_demux_002:src2_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	wire  [105:0] cmd_xbar_demux_002_src2_data;                                                                     // cmd_xbar_demux_002:src2_data -> cmd_xbar_mux_002:sink1_data
	wire    [4:0] cmd_xbar_demux_002_src2_channel;                                                                  // cmd_xbar_demux_002:src2_channel -> cmd_xbar_mux_002:sink1_channel
	wire          cmd_xbar_demux_002_src2_ready;                                                                    // cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_002:src2_ready
	wire          cmd_xbar_demux_002_src3_endofpacket;                                                              // cmd_xbar_demux_002:src3_endofpacket -> cmd_xbar_mux_003:sink2_endofpacket
	wire          cmd_xbar_demux_002_src3_valid;                                                                    // cmd_xbar_demux_002:src3_valid -> cmd_xbar_mux_003:sink2_valid
	wire          cmd_xbar_demux_002_src3_startofpacket;                                                            // cmd_xbar_demux_002:src3_startofpacket -> cmd_xbar_mux_003:sink2_startofpacket
	wire  [105:0] cmd_xbar_demux_002_src3_data;                                                                     // cmd_xbar_demux_002:src3_data -> cmd_xbar_mux_003:sink2_data
	wire    [4:0] cmd_xbar_demux_002_src3_channel;                                                                  // cmd_xbar_demux_002:src3_channel -> cmd_xbar_mux_003:sink2_channel
	wire          cmd_xbar_demux_002_src3_ready;                                                                    // cmd_xbar_mux_003:sink2_ready -> cmd_xbar_demux_002:src3_ready
	wire          cmd_xbar_demux_003_src0_endofpacket;                                                              // cmd_xbar_demux_003:src0_endofpacket -> cmd_xbar_mux_001:sink3_endofpacket
	wire          cmd_xbar_demux_003_src0_valid;                                                                    // cmd_xbar_demux_003:src0_valid -> cmd_xbar_mux_001:sink3_valid
	wire          cmd_xbar_demux_003_src0_startofpacket;                                                            // cmd_xbar_demux_003:src0_startofpacket -> cmd_xbar_mux_001:sink3_startofpacket
	wire  [105:0] cmd_xbar_demux_003_src0_data;                                                                     // cmd_xbar_demux_003:src0_data -> cmd_xbar_mux_001:sink3_data
	wire    [4:0] cmd_xbar_demux_003_src0_channel;                                                                  // cmd_xbar_demux_003:src0_channel -> cmd_xbar_mux_001:sink3_channel
	wire          cmd_xbar_demux_003_src0_ready;                                                                    // cmd_xbar_mux_001:sink3_ready -> cmd_xbar_demux_003:src0_ready
	wire          cmd_xbar_demux_003_src1_endofpacket;                                                              // cmd_xbar_demux_003:src1_endofpacket -> cmd_xbar_mux_003:sink3_endofpacket
	wire          cmd_xbar_demux_003_src1_valid;                                                                    // cmd_xbar_demux_003:src1_valid -> cmd_xbar_mux_003:sink3_valid
	wire          cmd_xbar_demux_003_src1_startofpacket;                                                            // cmd_xbar_demux_003:src1_startofpacket -> cmd_xbar_mux_003:sink3_startofpacket
	wire  [105:0] cmd_xbar_demux_003_src1_data;                                                                     // cmd_xbar_demux_003:src1_data -> cmd_xbar_mux_003:sink3_data
	wire    [4:0] cmd_xbar_demux_003_src1_channel;                                                                  // cmd_xbar_demux_003:src1_channel -> cmd_xbar_mux_003:sink3_channel
	wire          cmd_xbar_demux_003_src1_ready;                                                                    // cmd_xbar_mux_003:sink3_ready -> cmd_xbar_demux_003:src1_ready
	wire          rsp_xbar_demux_src0_endofpacket;                                                                  // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                        // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                                // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [105:0] rsp_xbar_demux_src0_data;                                                                         // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire    [4:0] rsp_xbar_demux_src0_channel;                                                                      // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire          rsp_xbar_demux_src0_ready;                                                                        // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire          rsp_xbar_demux_src1_endofpacket;                                                                  // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_002:sink0_endofpacket
	wire          rsp_xbar_demux_src1_valid;                                                                        // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_002:sink0_valid
	wire          rsp_xbar_demux_src1_startofpacket;                                                                // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_002:sink0_startofpacket
	wire  [105:0] rsp_xbar_demux_src1_data;                                                                         // rsp_xbar_demux:src1_data -> rsp_xbar_mux_002:sink0_data
	wire    [4:0] rsp_xbar_demux_src1_channel;                                                                      // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_002:sink0_channel
	wire          rsp_xbar_demux_src1_ready;                                                                        // rsp_xbar_mux_002:sink0_ready -> rsp_xbar_demux:src1_ready
	wire          rsp_xbar_demux_001_src0_endofpacket;                                                              // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                                    // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                                            // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [105:0] rsp_xbar_demux_001_src0_data;                                                                     // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire    [4:0] rsp_xbar_demux_001_src0_channel;                                                                  // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                                    // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire          rsp_xbar_demux_001_src1_endofpacket;                                                              // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire          rsp_xbar_demux_001_src1_valid;                                                                    // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire          rsp_xbar_demux_001_src1_startofpacket;                                                            // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [105:0] rsp_xbar_demux_001_src1_data;                                                                     // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink0_data
	wire    [4:0] rsp_xbar_demux_001_src1_channel;                                                                  // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire          rsp_xbar_demux_001_src1_ready;                                                                    // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux_001:src1_ready
	wire          rsp_xbar_demux_001_src2_endofpacket;                                                              // rsp_xbar_demux_001:src2_endofpacket -> rsp_xbar_mux_002:sink1_endofpacket
	wire          rsp_xbar_demux_001_src2_valid;                                                                    // rsp_xbar_demux_001:src2_valid -> rsp_xbar_mux_002:sink1_valid
	wire          rsp_xbar_demux_001_src2_startofpacket;                                                            // rsp_xbar_demux_001:src2_startofpacket -> rsp_xbar_mux_002:sink1_startofpacket
	wire  [105:0] rsp_xbar_demux_001_src2_data;                                                                     // rsp_xbar_demux_001:src2_data -> rsp_xbar_mux_002:sink1_data
	wire    [4:0] rsp_xbar_demux_001_src2_channel;                                                                  // rsp_xbar_demux_001:src2_channel -> rsp_xbar_mux_002:sink1_channel
	wire          rsp_xbar_demux_001_src2_ready;                                                                    // rsp_xbar_mux_002:sink1_ready -> rsp_xbar_demux_001:src2_ready
	wire          rsp_xbar_demux_001_src3_endofpacket;                                                              // rsp_xbar_demux_001:src3_endofpacket -> rsp_xbar_mux_003:sink0_endofpacket
	wire          rsp_xbar_demux_001_src3_valid;                                                                    // rsp_xbar_demux_001:src3_valid -> rsp_xbar_mux_003:sink0_valid
	wire          rsp_xbar_demux_001_src3_startofpacket;                                                            // rsp_xbar_demux_001:src3_startofpacket -> rsp_xbar_mux_003:sink0_startofpacket
	wire  [105:0] rsp_xbar_demux_001_src3_data;                                                                     // rsp_xbar_demux_001:src3_data -> rsp_xbar_mux_003:sink0_data
	wire    [4:0] rsp_xbar_demux_001_src3_channel;                                                                  // rsp_xbar_demux_001:src3_channel -> rsp_xbar_mux_003:sink0_channel
	wire          rsp_xbar_demux_001_src3_ready;                                                                    // rsp_xbar_mux_003:sink0_ready -> rsp_xbar_demux_001:src3_ready
	wire          rsp_xbar_demux_002_src0_endofpacket;                                                              // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire          rsp_xbar_demux_002_src0_valid;                                                                    // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire          rsp_xbar_demux_002_src0_startofpacket;                                                            // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [105:0] rsp_xbar_demux_002_src0_data;                                                                     // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire    [4:0] rsp_xbar_demux_002_src0_channel;                                                                  // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire          rsp_xbar_demux_002_src0_ready;                                                                    // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire          rsp_xbar_demux_002_src1_endofpacket;                                                              // rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_002:sink2_endofpacket
	wire          rsp_xbar_demux_002_src1_valid;                                                                    // rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_002:sink2_valid
	wire          rsp_xbar_demux_002_src1_startofpacket;                                                            // rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_002:sink2_startofpacket
	wire  [105:0] rsp_xbar_demux_002_src1_data;                                                                     // rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_002:sink2_data
	wire    [4:0] rsp_xbar_demux_002_src1_channel;                                                                  // rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_002:sink2_channel
	wire          rsp_xbar_demux_002_src1_ready;                                                                    // rsp_xbar_mux_002:sink2_ready -> rsp_xbar_demux_002:src1_ready
	wire          rsp_xbar_demux_003_src0_endofpacket;                                                              // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	wire          rsp_xbar_demux_003_src0_valid;                                                                    // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	wire          rsp_xbar_demux_003_src0_startofpacket;                                                            // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	wire  [105:0] rsp_xbar_demux_003_src0_data;                                                                     // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	wire    [4:0] rsp_xbar_demux_003_src0_channel;                                                                  // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	wire          rsp_xbar_demux_003_src0_ready;                                                                    // rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire          rsp_xbar_demux_003_src1_endofpacket;                                                              // rsp_xbar_demux_003:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire          rsp_xbar_demux_003_src1_valid;                                                                    // rsp_xbar_demux_003:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire          rsp_xbar_demux_003_src1_startofpacket;                                                            // rsp_xbar_demux_003:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [105:0] rsp_xbar_demux_003_src1_data;                                                                     // rsp_xbar_demux_003:src1_data -> rsp_xbar_mux_001:sink1_data
	wire    [4:0] rsp_xbar_demux_003_src1_channel;                                                                  // rsp_xbar_demux_003:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire          rsp_xbar_demux_003_src1_ready;                                                                    // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_003:src1_ready
	wire          rsp_xbar_demux_003_src2_endofpacket;                                                              // rsp_xbar_demux_003:src2_endofpacket -> rsp_xbar_mux_002:sink3_endofpacket
	wire          rsp_xbar_demux_003_src2_valid;                                                                    // rsp_xbar_demux_003:src2_valid -> rsp_xbar_mux_002:sink3_valid
	wire          rsp_xbar_demux_003_src2_startofpacket;                                                            // rsp_xbar_demux_003:src2_startofpacket -> rsp_xbar_mux_002:sink3_startofpacket
	wire  [105:0] rsp_xbar_demux_003_src2_data;                                                                     // rsp_xbar_demux_003:src2_data -> rsp_xbar_mux_002:sink3_data
	wire    [4:0] rsp_xbar_demux_003_src2_channel;                                                                  // rsp_xbar_demux_003:src2_channel -> rsp_xbar_mux_002:sink3_channel
	wire          rsp_xbar_demux_003_src2_ready;                                                                    // rsp_xbar_mux_002:sink3_ready -> rsp_xbar_demux_003:src2_ready
	wire          rsp_xbar_demux_003_src3_endofpacket;                                                              // rsp_xbar_demux_003:src3_endofpacket -> rsp_xbar_mux_003:sink1_endofpacket
	wire          rsp_xbar_demux_003_src3_valid;                                                                    // rsp_xbar_demux_003:src3_valid -> rsp_xbar_mux_003:sink1_valid
	wire          rsp_xbar_demux_003_src3_startofpacket;                                                            // rsp_xbar_demux_003:src3_startofpacket -> rsp_xbar_mux_003:sink1_startofpacket
	wire  [105:0] rsp_xbar_demux_003_src3_data;                                                                     // rsp_xbar_demux_003:src3_data -> rsp_xbar_mux_003:sink1_data
	wire    [4:0] rsp_xbar_demux_003_src3_channel;                                                                  // rsp_xbar_demux_003:src3_channel -> rsp_xbar_mux_003:sink1_channel
	wire          rsp_xbar_demux_003_src3_ready;                                                                    // rsp_xbar_mux_003:sink1_ready -> rsp_xbar_demux_003:src3_ready
	wire          addr_router_src_endofpacket;                                                                      // addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          addr_router_src_valid;                                                                            // addr_router:src_valid -> cmd_xbar_demux:sink_valid
	wire          addr_router_src_startofpacket;                                                                    // addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [105:0] addr_router_src_data;                                                                             // addr_router:src_data -> cmd_xbar_demux:sink_data
	wire    [4:0] addr_router_src_channel;                                                                          // addr_router:src_channel -> cmd_xbar_demux:sink_channel
	wire          addr_router_src_ready;                                                                            // cmd_xbar_demux:sink_ready -> addr_router:src_ready
	wire          rsp_xbar_mux_src_endofpacket;                                                                     // rsp_xbar_mux:src_endofpacket -> nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_src_valid;                                                                           // rsp_xbar_mux:src_valid -> nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_src_startofpacket;                                                                   // rsp_xbar_mux:src_startofpacket -> nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [105:0] rsp_xbar_mux_src_data;                                                                            // rsp_xbar_mux:src_data -> nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [4:0] rsp_xbar_mux_src_channel;                                                                         // rsp_xbar_mux:src_channel -> nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_src_ready;                                                                           // nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux:src_ready
	wire          addr_router_001_src_endofpacket;                                                                  // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          addr_router_001_src_valid;                                                                        // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire          addr_router_001_src_startofpacket;                                                                // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [105:0] addr_router_001_src_data;                                                                         // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire    [4:0] addr_router_001_src_channel;                                                                      // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire          addr_router_001_src_ready;                                                                        // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire          rsp_xbar_mux_001_src_endofpacket;                                                                 // rsp_xbar_mux_001:src_endofpacket -> dma_write_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_001_src_valid;                                                                       // rsp_xbar_mux_001:src_valid -> dma_write_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_001_src_startofpacket;                                                               // rsp_xbar_mux_001:src_startofpacket -> dma_write_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [105:0] rsp_xbar_mux_001_src_data;                                                                        // rsp_xbar_mux_001:src_data -> dma_write_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [4:0] rsp_xbar_mux_001_src_channel;                                                                     // rsp_xbar_mux_001:src_channel -> dma_write_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_001_src_ready;                                                                       // dma_write_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	wire          addr_router_002_src_endofpacket;                                                                  // addr_router_002:src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	wire          addr_router_002_src_valid;                                                                        // addr_router_002:src_valid -> cmd_xbar_demux_002:sink_valid
	wire          addr_router_002_src_startofpacket;                                                                // addr_router_002:src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	wire  [105:0] addr_router_002_src_data;                                                                         // addr_router_002:src_data -> cmd_xbar_demux_002:sink_data
	wire    [4:0] addr_router_002_src_channel;                                                                      // addr_router_002:src_channel -> cmd_xbar_demux_002:sink_channel
	wire          addr_router_002_src_ready;                                                                        // cmd_xbar_demux_002:sink_ready -> addr_router_002:src_ready
	wire          rsp_xbar_mux_002_src_endofpacket;                                                                 // rsp_xbar_mux_002:src_endofpacket -> nios2cpu_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_002_src_valid;                                                                       // rsp_xbar_mux_002:src_valid -> nios2cpu_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_002_src_startofpacket;                                                               // rsp_xbar_mux_002:src_startofpacket -> nios2cpu_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [105:0] rsp_xbar_mux_002_src_data;                                                                        // rsp_xbar_mux_002:src_data -> nios2cpu_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [4:0] rsp_xbar_mux_002_src_channel;                                                                     // rsp_xbar_mux_002:src_channel -> nios2cpu_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_002_src_ready;                                                                       // nios2cpu_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_002:src_ready
	wire          limiter_cmd_src_endofpacket;                                                                      // limiter:cmd_src_endofpacket -> cmd_xbar_demux_003:sink_endofpacket
	wire          limiter_cmd_src_startofpacket;                                                                    // limiter:cmd_src_startofpacket -> cmd_xbar_demux_003:sink_startofpacket
	wire  [105:0] limiter_cmd_src_data;                                                                             // limiter:cmd_src_data -> cmd_xbar_demux_003:sink_data
	wire    [4:0] limiter_cmd_src_channel;                                                                          // limiter:cmd_src_channel -> cmd_xbar_demux_003:sink_channel
	wire          limiter_cmd_src_ready;                                                                            // cmd_xbar_demux_003:sink_ready -> limiter:cmd_src_ready
	wire          rsp_xbar_mux_003_src_endofpacket;                                                                 // rsp_xbar_mux_003:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire          rsp_xbar_mux_003_src_valid;                                                                       // rsp_xbar_mux_003:src_valid -> limiter:rsp_sink_valid
	wire          rsp_xbar_mux_003_src_startofpacket;                                                               // rsp_xbar_mux_003:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [105:0] rsp_xbar_mux_003_src_data;                                                                        // rsp_xbar_mux_003:src_data -> limiter:rsp_sink_data
	wire    [4:0] rsp_xbar_mux_003_src_channel;                                                                     // rsp_xbar_mux_003:src_channel -> limiter:rsp_sink_channel
	wire          rsp_xbar_mux_003_src_ready;                                                                       // limiter:rsp_sink_ready -> rsp_xbar_mux_003:src_ready
	wire          cmd_xbar_mux_src_endofpacket;                                                                     // cmd_xbar_mux:src_endofpacket -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_src_valid;                                                                           // cmd_xbar_mux:src_valid -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_src_startofpacket;                                                                   // cmd_xbar_mux:src_startofpacket -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [105:0] cmd_xbar_mux_src_data;                                                                            // cmd_xbar_mux:src_data -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire    [4:0] cmd_xbar_mux_src_channel;                                                                         // cmd_xbar_mux:src_channel -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_src_ready;                                                                           // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire          id_router_src_endofpacket;                                                                        // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          id_router_src_valid;                                                                              // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire          id_router_src_startofpacket;                                                                      // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [105:0] id_router_src_data;                                                                               // id_router:src_data -> rsp_xbar_demux:sink_data
	wire    [4:0] id_router_src_channel;                                                                            // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire          id_router_src_ready;                                                                              // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire          cmd_xbar_mux_002_src_endofpacket;                                                                 // cmd_xbar_mux_002:src_endofpacket -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_002_src_valid;                                                                       // cmd_xbar_mux_002:src_valid -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_002_src_startofpacket;                                                               // cmd_xbar_mux_002:src_startofpacket -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [105:0] cmd_xbar_mux_002_src_data;                                                                        // cmd_xbar_mux_002:src_data -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire    [4:0] cmd_xbar_mux_002_src_channel;                                                                     // cmd_xbar_mux_002:src_channel -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_002_src_ready;                                                                       // dma_control_port_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_002:src_ready
	wire          id_router_002_src_endofpacket;                                                                    // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire          id_router_002_src_valid;                                                                          // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire          id_router_002_src_startofpacket;                                                                  // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [105:0] id_router_002_src_data;                                                                           // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire    [4:0] id_router_002_src_channel;                                                                        // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire          id_router_002_src_ready;                                                                          // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire          cmd_xbar_mux_003_src_endofpacket;                                                                 // cmd_xbar_mux_003:src_endofpacket -> burst_adapter_001:sink0_endofpacket
	wire          cmd_xbar_mux_003_src_valid;                                                                       // cmd_xbar_mux_003:src_valid -> burst_adapter_001:sink0_valid
	wire          cmd_xbar_mux_003_src_startofpacket;                                                               // cmd_xbar_mux_003:src_startofpacket -> burst_adapter_001:sink0_startofpacket
	wire  [105:0] cmd_xbar_mux_003_src_data;                                                                        // cmd_xbar_mux_003:src_data -> burst_adapter_001:sink0_data
	wire    [4:0] cmd_xbar_mux_003_src_channel;                                                                     // cmd_xbar_mux_003:src_channel -> burst_adapter_001:sink0_channel
	wire          cmd_xbar_mux_003_src_ready;                                                                       // burst_adapter_001:sink0_ready -> cmd_xbar_mux_003:src_ready
	wire          id_router_003_src_endofpacket;                                                                    // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire          id_router_003_src_valid;                                                                          // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire          id_router_003_src_startofpacket;                                                                  // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [105:0] id_router_003_src_data;                                                                           // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire    [4:0] id_router_003_src_channel;                                                                        // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire          id_router_003_src_ready;                                                                          // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire          crosser_out_ready;                                                                                // syspll_pll_slave_translator_avalon_universal_slave_0_agent:cp_ready -> crosser:out_ready
	wire          id_router_004_src_endofpacket;                                                                    // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire          id_router_004_src_valid;                                                                          // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire          id_router_004_src_startofpacket;                                                                  // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [105:0] id_router_004_src_data;                                                                           // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire    [4:0] id_router_004_src_channel;                                                                        // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire          id_router_004_src_ready;                                                                          // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire          cmd_xbar_demux_004_src0_endofpacket;                                                              // cmd_xbar_demux_004:src0_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_004_src0_valid;                                                                    // cmd_xbar_demux_004:src0_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_004_src0_startofpacket;                                                            // cmd_xbar_demux_004:src0_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [82:0] cmd_xbar_demux_004_src0_data;                                                                     // cmd_xbar_demux_004:src0_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [10:0] cmd_xbar_demux_004_src0_channel;                                                                  // cmd_xbar_demux_004:src0_channel -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_004_src1_endofpacket;                                                              // cmd_xbar_demux_004:src1_endofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_004_src1_valid;                                                                    // cmd_xbar_demux_004:src1_valid -> timer_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_004_src1_startofpacket;                                                            // cmd_xbar_demux_004:src1_startofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [82:0] cmd_xbar_demux_004_src1_data;                                                                     // cmd_xbar_demux_004:src1_data -> timer_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [10:0] cmd_xbar_demux_004_src1_channel;                                                                  // cmd_xbar_demux_004:src1_channel -> timer_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_004_src2_endofpacket;                                                              // cmd_xbar_demux_004:src2_endofpacket -> uart0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_004_src2_valid;                                                                    // cmd_xbar_demux_004:src2_valid -> uart0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_004_src2_startofpacket;                                                            // cmd_xbar_demux_004:src2_startofpacket -> uart0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [82:0] cmd_xbar_demux_004_src2_data;                                                                     // cmd_xbar_demux_004:src2_data -> uart0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [10:0] cmd_xbar_demux_004_src2_channel;                                                                  // cmd_xbar_demux_004:src2_channel -> uart0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_004_src3_endofpacket;                                                              // cmd_xbar_demux_004:src3_endofpacket -> sw_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_004_src3_valid;                                                                    // cmd_xbar_demux_004:src3_valid -> sw_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_004_src3_startofpacket;                                                            // cmd_xbar_demux_004:src3_startofpacket -> sw_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [82:0] cmd_xbar_demux_004_src3_data;                                                                     // cmd_xbar_demux_004:src3_data -> sw_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [10:0] cmd_xbar_demux_004_src3_channel;                                                                  // cmd_xbar_demux_004:src3_channel -> sw_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_004_src4_endofpacket;                                                              // cmd_xbar_demux_004:src4_endofpacket -> led_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_004_src4_valid;                                                                    // cmd_xbar_demux_004:src4_valid -> led_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_004_src4_startofpacket;                                                            // cmd_xbar_demux_004:src4_startofpacket -> led_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [82:0] cmd_xbar_demux_004_src4_data;                                                                     // cmd_xbar_demux_004:src4_data -> led_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [10:0] cmd_xbar_demux_004_src4_channel;                                                                  // cmd_xbar_demux_004:src4_channel -> led_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_004_src5_endofpacket;                                                              // cmd_xbar_demux_004:src5_endofpacket -> button1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_004_src5_valid;                                                                    // cmd_xbar_demux_004:src5_valid -> button1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_004_src5_startofpacket;                                                            // cmd_xbar_demux_004:src5_startofpacket -> button1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [82:0] cmd_xbar_demux_004_src5_data;                                                                     // cmd_xbar_demux_004:src5_data -> button1_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [10:0] cmd_xbar_demux_004_src5_channel;                                                                  // cmd_xbar_demux_004:src5_channel -> button1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_004_src6_endofpacket;                                                              // cmd_xbar_demux_004:src6_endofpacket -> button2_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_004_src6_valid;                                                                    // cmd_xbar_demux_004:src6_valid -> button2_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_004_src6_startofpacket;                                                            // cmd_xbar_demux_004:src6_startofpacket -> button2_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [82:0] cmd_xbar_demux_004_src6_data;                                                                     // cmd_xbar_demux_004:src6_data -> button2_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [10:0] cmd_xbar_demux_004_src6_channel;                                                                  // cmd_xbar_demux_004:src6_channel -> button2_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_004_src7_endofpacket;                                                              // cmd_xbar_demux_004:src7_endofpacket -> hex0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_004_src7_valid;                                                                    // cmd_xbar_demux_004:src7_valid -> hex0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_004_src7_startofpacket;                                                            // cmd_xbar_demux_004:src7_startofpacket -> hex0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [82:0] cmd_xbar_demux_004_src7_data;                                                                     // cmd_xbar_demux_004:src7_data -> hex0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [10:0] cmd_xbar_demux_004_src7_channel;                                                                  // cmd_xbar_demux_004:src7_channel -> hex0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_004_src8_endofpacket;                                                              // cmd_xbar_demux_004:src8_endofpacket -> hex1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_004_src8_valid;                                                                    // cmd_xbar_demux_004:src8_valid -> hex1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_004_src8_startofpacket;                                                            // cmd_xbar_demux_004:src8_startofpacket -> hex1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [82:0] cmd_xbar_demux_004_src8_data;                                                                     // cmd_xbar_demux_004:src8_data -> hex1_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [10:0] cmd_xbar_demux_004_src8_channel;                                                                  // cmd_xbar_demux_004:src8_channel -> hex1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_004_src9_endofpacket;                                                              // cmd_xbar_demux_004:src9_endofpacket -> hex2_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_004_src9_valid;                                                                    // cmd_xbar_demux_004:src9_valid -> hex2_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_004_src9_startofpacket;                                                            // cmd_xbar_demux_004:src9_startofpacket -> hex2_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [82:0] cmd_xbar_demux_004_src9_data;                                                                     // cmd_xbar_demux_004:src9_data -> hex2_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [10:0] cmd_xbar_demux_004_src9_channel;                                                                  // cmd_xbar_demux_004:src9_channel -> hex2_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_004_src10_endofpacket;                                                             // cmd_xbar_demux_004:src10_endofpacket -> hex3_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_004_src10_valid;                                                                   // cmd_xbar_demux_004:src10_valid -> hex3_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_004_src10_startofpacket;                                                           // cmd_xbar_demux_004:src10_startofpacket -> hex3_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [82:0] cmd_xbar_demux_004_src10_data;                                                                    // cmd_xbar_demux_004:src10_data -> hex3_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [10:0] cmd_xbar_demux_004_src10_channel;                                                                 // cmd_xbar_demux_004:src10_channel -> hex3_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rsp_xbar_demux_005_src0_endofpacket;                                                              // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_004:sink0_endofpacket
	wire          rsp_xbar_demux_005_src0_valid;                                                                    // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_004:sink0_valid
	wire          rsp_xbar_demux_005_src0_startofpacket;                                                            // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_004:sink0_startofpacket
	wire   [82:0] rsp_xbar_demux_005_src0_data;                                                                     // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_004:sink0_data
	wire   [10:0] rsp_xbar_demux_005_src0_channel;                                                                  // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_004:sink0_channel
	wire          rsp_xbar_demux_005_src0_ready;                                                                    // rsp_xbar_mux_004:sink0_ready -> rsp_xbar_demux_005:src0_ready
	wire          rsp_xbar_demux_006_src0_endofpacket;                                                              // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_004:sink1_endofpacket
	wire          rsp_xbar_demux_006_src0_valid;                                                                    // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_004:sink1_valid
	wire          rsp_xbar_demux_006_src0_startofpacket;                                                            // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_004:sink1_startofpacket
	wire   [82:0] rsp_xbar_demux_006_src0_data;                                                                     // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_004:sink1_data
	wire   [10:0] rsp_xbar_demux_006_src0_channel;                                                                  // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_004:sink1_channel
	wire          rsp_xbar_demux_006_src0_ready;                                                                    // rsp_xbar_mux_004:sink1_ready -> rsp_xbar_demux_006:src0_ready
	wire          rsp_xbar_demux_007_src0_endofpacket;                                                              // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_004:sink2_endofpacket
	wire          rsp_xbar_demux_007_src0_valid;                                                                    // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_004:sink2_valid
	wire          rsp_xbar_demux_007_src0_startofpacket;                                                            // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_004:sink2_startofpacket
	wire   [82:0] rsp_xbar_demux_007_src0_data;                                                                     // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_004:sink2_data
	wire   [10:0] rsp_xbar_demux_007_src0_channel;                                                                  // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_004:sink2_channel
	wire          rsp_xbar_demux_007_src0_ready;                                                                    // rsp_xbar_mux_004:sink2_ready -> rsp_xbar_demux_007:src0_ready
	wire          rsp_xbar_demux_008_src0_endofpacket;                                                              // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_004:sink3_endofpacket
	wire          rsp_xbar_demux_008_src0_valid;                                                                    // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_004:sink3_valid
	wire          rsp_xbar_demux_008_src0_startofpacket;                                                            // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_004:sink3_startofpacket
	wire   [82:0] rsp_xbar_demux_008_src0_data;                                                                     // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_004:sink3_data
	wire   [10:0] rsp_xbar_demux_008_src0_channel;                                                                  // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_004:sink3_channel
	wire          rsp_xbar_demux_008_src0_ready;                                                                    // rsp_xbar_mux_004:sink3_ready -> rsp_xbar_demux_008:src0_ready
	wire          rsp_xbar_demux_009_src0_endofpacket;                                                              // rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_004:sink4_endofpacket
	wire          rsp_xbar_demux_009_src0_valid;                                                                    // rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_004:sink4_valid
	wire          rsp_xbar_demux_009_src0_startofpacket;                                                            // rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_004:sink4_startofpacket
	wire   [82:0] rsp_xbar_demux_009_src0_data;                                                                     // rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_004:sink4_data
	wire   [10:0] rsp_xbar_demux_009_src0_channel;                                                                  // rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_004:sink4_channel
	wire          rsp_xbar_demux_009_src0_ready;                                                                    // rsp_xbar_mux_004:sink4_ready -> rsp_xbar_demux_009:src0_ready
	wire          rsp_xbar_demux_010_src0_endofpacket;                                                              // rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux_004:sink5_endofpacket
	wire          rsp_xbar_demux_010_src0_valid;                                                                    // rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux_004:sink5_valid
	wire          rsp_xbar_demux_010_src0_startofpacket;                                                            // rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux_004:sink5_startofpacket
	wire   [82:0] rsp_xbar_demux_010_src0_data;                                                                     // rsp_xbar_demux_010:src0_data -> rsp_xbar_mux_004:sink5_data
	wire   [10:0] rsp_xbar_demux_010_src0_channel;                                                                  // rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux_004:sink5_channel
	wire          rsp_xbar_demux_010_src0_ready;                                                                    // rsp_xbar_mux_004:sink5_ready -> rsp_xbar_demux_010:src0_ready
	wire          rsp_xbar_demux_011_src0_endofpacket;                                                              // rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux_004:sink6_endofpacket
	wire          rsp_xbar_demux_011_src0_valid;                                                                    // rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux_004:sink6_valid
	wire          rsp_xbar_demux_011_src0_startofpacket;                                                            // rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux_004:sink6_startofpacket
	wire   [82:0] rsp_xbar_demux_011_src0_data;                                                                     // rsp_xbar_demux_011:src0_data -> rsp_xbar_mux_004:sink6_data
	wire   [10:0] rsp_xbar_demux_011_src0_channel;                                                                  // rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux_004:sink6_channel
	wire          rsp_xbar_demux_011_src0_ready;                                                                    // rsp_xbar_mux_004:sink6_ready -> rsp_xbar_demux_011:src0_ready
	wire          rsp_xbar_demux_012_src0_endofpacket;                                                              // rsp_xbar_demux_012:src0_endofpacket -> rsp_xbar_mux_004:sink7_endofpacket
	wire          rsp_xbar_demux_012_src0_valid;                                                                    // rsp_xbar_demux_012:src0_valid -> rsp_xbar_mux_004:sink7_valid
	wire          rsp_xbar_demux_012_src0_startofpacket;                                                            // rsp_xbar_demux_012:src0_startofpacket -> rsp_xbar_mux_004:sink7_startofpacket
	wire   [82:0] rsp_xbar_demux_012_src0_data;                                                                     // rsp_xbar_demux_012:src0_data -> rsp_xbar_mux_004:sink7_data
	wire   [10:0] rsp_xbar_demux_012_src0_channel;                                                                  // rsp_xbar_demux_012:src0_channel -> rsp_xbar_mux_004:sink7_channel
	wire          rsp_xbar_demux_012_src0_ready;                                                                    // rsp_xbar_mux_004:sink7_ready -> rsp_xbar_demux_012:src0_ready
	wire          rsp_xbar_demux_013_src0_endofpacket;                                                              // rsp_xbar_demux_013:src0_endofpacket -> rsp_xbar_mux_004:sink8_endofpacket
	wire          rsp_xbar_demux_013_src0_valid;                                                                    // rsp_xbar_demux_013:src0_valid -> rsp_xbar_mux_004:sink8_valid
	wire          rsp_xbar_demux_013_src0_startofpacket;                                                            // rsp_xbar_demux_013:src0_startofpacket -> rsp_xbar_mux_004:sink8_startofpacket
	wire   [82:0] rsp_xbar_demux_013_src0_data;                                                                     // rsp_xbar_demux_013:src0_data -> rsp_xbar_mux_004:sink8_data
	wire   [10:0] rsp_xbar_demux_013_src0_channel;                                                                  // rsp_xbar_demux_013:src0_channel -> rsp_xbar_mux_004:sink8_channel
	wire          rsp_xbar_demux_013_src0_ready;                                                                    // rsp_xbar_mux_004:sink8_ready -> rsp_xbar_demux_013:src0_ready
	wire          rsp_xbar_demux_014_src0_endofpacket;                                                              // rsp_xbar_demux_014:src0_endofpacket -> rsp_xbar_mux_004:sink9_endofpacket
	wire          rsp_xbar_demux_014_src0_valid;                                                                    // rsp_xbar_demux_014:src0_valid -> rsp_xbar_mux_004:sink9_valid
	wire          rsp_xbar_demux_014_src0_startofpacket;                                                            // rsp_xbar_demux_014:src0_startofpacket -> rsp_xbar_mux_004:sink9_startofpacket
	wire   [82:0] rsp_xbar_demux_014_src0_data;                                                                     // rsp_xbar_demux_014:src0_data -> rsp_xbar_mux_004:sink9_data
	wire   [10:0] rsp_xbar_demux_014_src0_channel;                                                                  // rsp_xbar_demux_014:src0_channel -> rsp_xbar_mux_004:sink9_channel
	wire          rsp_xbar_demux_014_src0_ready;                                                                    // rsp_xbar_mux_004:sink9_ready -> rsp_xbar_demux_014:src0_ready
	wire          rsp_xbar_demux_015_src0_endofpacket;                                                              // rsp_xbar_demux_015:src0_endofpacket -> rsp_xbar_mux_004:sink10_endofpacket
	wire          rsp_xbar_demux_015_src0_valid;                                                                    // rsp_xbar_demux_015:src0_valid -> rsp_xbar_mux_004:sink10_valid
	wire          rsp_xbar_demux_015_src0_startofpacket;                                                            // rsp_xbar_demux_015:src0_startofpacket -> rsp_xbar_mux_004:sink10_startofpacket
	wire   [82:0] rsp_xbar_demux_015_src0_data;                                                                     // rsp_xbar_demux_015:src0_data -> rsp_xbar_mux_004:sink10_data
	wire   [10:0] rsp_xbar_demux_015_src0_channel;                                                                  // rsp_xbar_demux_015:src0_channel -> rsp_xbar_mux_004:sink10_channel
	wire          rsp_xbar_demux_015_src0_ready;                                                                    // rsp_xbar_mux_004:sink10_ready -> rsp_xbar_demux_015:src0_ready
	wire          limiter_001_cmd_src_endofpacket;                                                                  // limiter_001:cmd_src_endofpacket -> cmd_xbar_demux_004:sink_endofpacket
	wire          limiter_001_cmd_src_startofpacket;                                                                // limiter_001:cmd_src_startofpacket -> cmd_xbar_demux_004:sink_startofpacket
	wire   [82:0] limiter_001_cmd_src_data;                                                                         // limiter_001:cmd_src_data -> cmd_xbar_demux_004:sink_data
	wire   [10:0] limiter_001_cmd_src_channel;                                                                      // limiter_001:cmd_src_channel -> cmd_xbar_demux_004:sink_channel
	wire          limiter_001_cmd_src_ready;                                                                        // cmd_xbar_demux_004:sink_ready -> limiter_001:cmd_src_ready
	wire          rsp_xbar_mux_004_src_endofpacket;                                                                 // rsp_xbar_mux_004:src_endofpacket -> limiter_001:rsp_sink_endofpacket
	wire          rsp_xbar_mux_004_src_valid;                                                                       // rsp_xbar_mux_004:src_valid -> limiter_001:rsp_sink_valid
	wire          rsp_xbar_mux_004_src_startofpacket;                                                               // rsp_xbar_mux_004:src_startofpacket -> limiter_001:rsp_sink_startofpacket
	wire   [82:0] rsp_xbar_mux_004_src_data;                                                                        // rsp_xbar_mux_004:src_data -> limiter_001:rsp_sink_data
	wire   [10:0] rsp_xbar_mux_004_src_channel;                                                                     // rsp_xbar_mux_004:src_channel -> limiter_001:rsp_sink_channel
	wire          rsp_xbar_mux_004_src_ready;                                                                       // limiter_001:rsp_sink_ready -> rsp_xbar_mux_004:src_ready
	wire          cmd_xbar_demux_004_src0_ready;                                                                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_004:src0_ready
	wire          id_router_005_src_endofpacket;                                                                    // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire          id_router_005_src_valid;                                                                          // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire          id_router_005_src_startofpacket;                                                                  // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire   [82:0] id_router_005_src_data;                                                                           // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire   [10:0] id_router_005_src_channel;                                                                        // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire          id_router_005_src_ready;                                                                          // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire          cmd_xbar_demux_004_src1_ready;                                                                    // timer_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_004:src1_ready
	wire          id_router_006_src_endofpacket;                                                                    // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire          id_router_006_src_valid;                                                                          // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire          id_router_006_src_startofpacket;                                                                  // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire   [82:0] id_router_006_src_data;                                                                           // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire   [10:0] id_router_006_src_channel;                                                                        // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire          id_router_006_src_ready;                                                                          // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire          cmd_xbar_demux_004_src2_ready;                                                                    // uart0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_004:src2_ready
	wire          id_router_007_src_endofpacket;                                                                    // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire          id_router_007_src_valid;                                                                          // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire          id_router_007_src_startofpacket;                                                                  // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire   [82:0] id_router_007_src_data;                                                                           // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire   [10:0] id_router_007_src_channel;                                                                        // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire          id_router_007_src_ready;                                                                          // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire          cmd_xbar_demux_004_src3_ready;                                                                    // sw_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_004:src3_ready
	wire          id_router_008_src_endofpacket;                                                                    // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire          id_router_008_src_valid;                                                                          // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire          id_router_008_src_startofpacket;                                                                  // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire   [82:0] id_router_008_src_data;                                                                           // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire   [10:0] id_router_008_src_channel;                                                                        // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire          id_router_008_src_ready;                                                                          // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire          cmd_xbar_demux_004_src4_ready;                                                                    // led_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_004:src4_ready
	wire          id_router_009_src_endofpacket;                                                                    // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire          id_router_009_src_valid;                                                                          // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire          id_router_009_src_startofpacket;                                                                  // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire   [82:0] id_router_009_src_data;                                                                           // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire   [10:0] id_router_009_src_channel;                                                                        // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire          id_router_009_src_ready;                                                                          // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire          cmd_xbar_demux_004_src5_ready;                                                                    // button1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_004:src5_ready
	wire          id_router_010_src_endofpacket;                                                                    // id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire          id_router_010_src_valid;                                                                          // id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	wire          id_router_010_src_startofpacket;                                                                  // id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire   [82:0] id_router_010_src_data;                                                                           // id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	wire   [10:0] id_router_010_src_channel;                                                                        // id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	wire          id_router_010_src_ready;                                                                          // rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	wire          cmd_xbar_demux_004_src6_ready;                                                                    // button2_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_004:src6_ready
	wire          id_router_011_src_endofpacket;                                                                    // id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	wire          id_router_011_src_valid;                                                                          // id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	wire          id_router_011_src_startofpacket;                                                                  // id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	wire   [82:0] id_router_011_src_data;                                                                           // id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	wire   [10:0] id_router_011_src_channel;                                                                        // id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	wire          id_router_011_src_ready;                                                                          // rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	wire          cmd_xbar_demux_004_src7_ready;                                                                    // hex0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_004:src7_ready
	wire          id_router_012_src_endofpacket;                                                                    // id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	wire          id_router_012_src_valid;                                                                          // id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	wire          id_router_012_src_startofpacket;                                                                  // id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	wire   [82:0] id_router_012_src_data;                                                                           // id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	wire   [10:0] id_router_012_src_channel;                                                                        // id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	wire          id_router_012_src_ready;                                                                          // rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	wire          cmd_xbar_demux_004_src8_ready;                                                                    // hex1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_004:src8_ready
	wire          id_router_013_src_endofpacket;                                                                    // id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	wire          id_router_013_src_valid;                                                                          // id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	wire          id_router_013_src_startofpacket;                                                                  // id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	wire   [82:0] id_router_013_src_data;                                                                           // id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	wire   [10:0] id_router_013_src_channel;                                                                        // id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	wire          id_router_013_src_ready;                                                                          // rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	wire          cmd_xbar_demux_004_src9_ready;                                                                    // hex2_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_004:src9_ready
	wire          id_router_014_src_endofpacket;                                                                    // id_router_014:src_endofpacket -> rsp_xbar_demux_014:sink_endofpacket
	wire          id_router_014_src_valid;                                                                          // id_router_014:src_valid -> rsp_xbar_demux_014:sink_valid
	wire          id_router_014_src_startofpacket;                                                                  // id_router_014:src_startofpacket -> rsp_xbar_demux_014:sink_startofpacket
	wire   [82:0] id_router_014_src_data;                                                                           // id_router_014:src_data -> rsp_xbar_demux_014:sink_data
	wire   [10:0] id_router_014_src_channel;                                                                        // id_router_014:src_channel -> rsp_xbar_demux_014:sink_channel
	wire          id_router_014_src_ready;                                                                          // rsp_xbar_demux_014:sink_ready -> id_router_014:src_ready
	wire          cmd_xbar_demux_004_src10_ready;                                                                   // hex3_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_004:src10_ready
	wire          id_router_015_src_endofpacket;                                                                    // id_router_015:src_endofpacket -> rsp_xbar_demux_015:sink_endofpacket
	wire          id_router_015_src_valid;                                                                          // id_router_015:src_valid -> rsp_xbar_demux_015:sink_valid
	wire          id_router_015_src_startofpacket;                                                                  // id_router_015:src_startofpacket -> rsp_xbar_demux_015:sink_startofpacket
	wire   [82:0] id_router_015_src_data;                                                                           // id_router_015:src_data -> rsp_xbar_demux_015:sink_data
	wire   [10:0] id_router_015_src_channel;                                                                        // id_router_015:src_channel -> rsp_xbar_demux_015:sink_channel
	wire          id_router_015_src_ready;                                                                          // rsp_xbar_demux_015:sink_ready -> id_router_015:src_ready
	wire          cmd_xbar_mux_001_src_endofpacket;                                                                 // cmd_xbar_mux_001:src_endofpacket -> width_adapter:in_endofpacket
	wire          cmd_xbar_mux_001_src_valid;                                                                       // cmd_xbar_mux_001:src_valid -> width_adapter:in_valid
	wire          cmd_xbar_mux_001_src_startofpacket;                                                               // cmd_xbar_mux_001:src_startofpacket -> width_adapter:in_startofpacket
	wire  [105:0] cmd_xbar_mux_001_src_data;                                                                        // cmd_xbar_mux_001:src_data -> width_adapter:in_data
	wire    [4:0] cmd_xbar_mux_001_src_channel;                                                                     // cmd_xbar_mux_001:src_channel -> width_adapter:in_channel
	wire          cmd_xbar_mux_001_src_ready;                                                                       // width_adapter:in_ready -> cmd_xbar_mux_001:src_ready
	wire          width_adapter_src_endofpacket;                                                                    // width_adapter:out_endofpacket -> burst_adapter:sink0_endofpacket
	wire          width_adapter_src_valid;                                                                          // width_adapter:out_valid -> burst_adapter:sink0_valid
	wire          width_adapter_src_startofpacket;                                                                  // width_adapter:out_startofpacket -> burst_adapter:sink0_startofpacket
	wire   [87:0] width_adapter_src_data;                                                                           // width_adapter:out_data -> burst_adapter:sink0_data
	wire          width_adapter_src_ready;                                                                          // burst_adapter:sink0_ready -> width_adapter:out_ready
	wire    [4:0] width_adapter_src_channel;                                                                        // width_adapter:out_channel -> burst_adapter:sink0_channel
	wire          id_router_001_src_endofpacket;                                                                    // id_router_001:src_endofpacket -> width_adapter_001:in_endofpacket
	wire          id_router_001_src_valid;                                                                          // id_router_001:src_valid -> width_adapter_001:in_valid
	wire          id_router_001_src_startofpacket;                                                                  // id_router_001:src_startofpacket -> width_adapter_001:in_startofpacket
	wire   [87:0] id_router_001_src_data;                                                                           // id_router_001:src_data -> width_adapter_001:in_data
	wire    [4:0] id_router_001_src_channel;                                                                        // id_router_001:src_channel -> width_adapter_001:in_channel
	wire          id_router_001_src_ready;                                                                          // width_adapter_001:in_ready -> id_router_001:src_ready
	wire          width_adapter_001_src_endofpacket;                                                                // width_adapter_001:out_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          width_adapter_001_src_valid;                                                                      // width_adapter_001:out_valid -> rsp_xbar_demux_001:sink_valid
	wire          width_adapter_001_src_startofpacket;                                                              // width_adapter_001:out_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [105:0] width_adapter_001_src_data;                                                                       // width_adapter_001:out_data -> rsp_xbar_demux_001:sink_data
	wire          width_adapter_001_src_ready;                                                                      // rsp_xbar_demux_001:sink_ready -> width_adapter_001:out_ready
	wire    [4:0] width_adapter_001_src_channel;                                                                    // width_adapter_001:out_channel -> rsp_xbar_demux_001:sink_channel
	wire          crosser_out_endofpacket;                                                                          // crosser:out_endofpacket -> syspll_pll_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_out_valid;                                                                                // crosser:out_valid -> syspll_pll_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_out_startofpacket;                                                                        // crosser:out_startofpacket -> syspll_pll_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [105:0] crosser_out_data;                                                                                 // crosser:out_data -> syspll_pll_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire    [4:0] crosser_out_channel;                                                                              // crosser:out_channel -> syspll_pll_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_002_src4_endofpacket;                                                              // cmd_xbar_demux_002:src4_endofpacket -> crosser:in_endofpacket
	wire          cmd_xbar_demux_002_src4_valid;                                                                    // cmd_xbar_demux_002:src4_valid -> crosser:in_valid
	wire          cmd_xbar_demux_002_src4_startofpacket;                                                            // cmd_xbar_demux_002:src4_startofpacket -> crosser:in_startofpacket
	wire  [105:0] cmd_xbar_demux_002_src4_data;                                                                     // cmd_xbar_demux_002:src4_data -> crosser:in_data
	wire    [4:0] cmd_xbar_demux_002_src4_channel;                                                                  // cmd_xbar_demux_002:src4_channel -> crosser:in_channel
	wire          cmd_xbar_demux_002_src4_ready;                                                                    // crosser:in_ready -> cmd_xbar_demux_002:src4_ready
	wire          crosser_001_out_endofpacket;                                                                      // crosser_001:out_endofpacket -> rsp_xbar_mux_002:sink4_endofpacket
	wire          crosser_001_out_valid;                                                                            // crosser_001:out_valid -> rsp_xbar_mux_002:sink4_valid
	wire          crosser_001_out_startofpacket;                                                                    // crosser_001:out_startofpacket -> rsp_xbar_mux_002:sink4_startofpacket
	wire  [105:0] crosser_001_out_data;                                                                             // crosser_001:out_data -> rsp_xbar_mux_002:sink4_data
	wire    [4:0] crosser_001_out_channel;                                                                          // crosser_001:out_channel -> rsp_xbar_mux_002:sink4_channel
	wire          crosser_001_out_ready;                                                                            // rsp_xbar_mux_002:sink4_ready -> crosser_001:out_ready
	wire          rsp_xbar_demux_004_src0_endofpacket;                                                              // rsp_xbar_demux_004:src0_endofpacket -> crosser_001:in_endofpacket
	wire          rsp_xbar_demux_004_src0_valid;                                                                    // rsp_xbar_demux_004:src0_valid -> crosser_001:in_valid
	wire          rsp_xbar_demux_004_src0_startofpacket;                                                            // rsp_xbar_demux_004:src0_startofpacket -> crosser_001:in_startofpacket
	wire  [105:0] rsp_xbar_demux_004_src0_data;                                                                     // rsp_xbar_demux_004:src0_data -> crosser_001:in_data
	wire    [4:0] rsp_xbar_demux_004_src0_channel;                                                                  // rsp_xbar_demux_004:src0_channel -> crosser_001:in_channel
	wire          rsp_xbar_demux_004_src0_ready;                                                                    // crosser_001:in_ready -> rsp_xbar_demux_004:src0_ready
	wire    [4:0] limiter_cmd_valid_data;                                                                           // limiter:cmd_src_valid -> cmd_xbar_demux_003:sink_valid
	wire   [10:0] limiter_001_cmd_valid_data;                                                                       // limiter_001:cmd_src_valid -> cmd_xbar_demux_004:sink_valid
	wire          irq_mapper_receiver0_irq;                                                                         // dma:dma_ctl_irq -> irq_mapper:receiver0_irq
	wire          irq_mapper_receiver1_irq;                                                                         // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire          irq_mapper_receiver2_irq;                                                                         // timer:irq -> irq_mapper:receiver2_irq
	wire          irq_mapper_receiver3_irq;                                                                         // uart0:irq -> irq_mapper:receiver3_irq
	wire          irq_mapper_receiver4_irq;                                                                         // button1:irq -> irq_mapper:receiver4_irq
	wire   [31:0] nios2cpu_d_irq_irq;                                                                               // irq_mapper:sender_irq -> nios2cpu:d_irq

	DE0Qsys_syspll syspll (
		.clk       (clk_50m_clk),                                               //       inclk_interface.clk
		.reset     (rst_controller_reset_out_reset),                            // inclk_interface_reset.reset
		.read      (syspll_pll_slave_translator_avalon_anti_slave_0_read),      //             pll_slave.read
		.write     (syspll_pll_slave_translator_avalon_anti_slave_0_write),     //                      .write
		.address   (syspll_pll_slave_translator_avalon_anti_slave_0_address),   //                      .address
		.readdata  (syspll_pll_slave_translator_avalon_anti_slave_0_readdata),  //                      .readdata
		.writedata (syspll_pll_slave_translator_avalon_anti_slave_0_writedata), //                      .writedata
		.c0        (syspll_c0_clk),                                             //                    c0.clk
		.c1        (dram_clk_clk),                                              //                    c1.clk
		.c2        (),                                                          //                    c2.clk
		.areset    (areset_export),                                             //        areset_conduit.export
		.locked    (locked_export),                                             //        locked_conduit.export
		.phasedone (phasedone_export)                                           //     phasedone_conduit.export
	);

	DE0Qsys_nios2cpu nios2cpu (
		.clk                                   (syspll_c0_clk),                                                         //                       clk.clk
		.reset_n                               (~rst_controller_001_reset_out_reset),                                   //                   reset_n.reset_n
		.d_address                             (nios2cpu_data_master_address),                                          //               data_master.address
		.d_byteenable                          (nios2cpu_data_master_byteenable),                                       //                          .byteenable
		.d_read                                (nios2cpu_data_master_read),                                             //                          .read
		.d_readdata                            (nios2cpu_data_master_readdata),                                         //                          .readdata
		.d_waitrequest                         (nios2cpu_data_master_waitrequest),                                      //                          .waitrequest
		.d_write                               (nios2cpu_data_master_write),                                            //                          .write
		.d_writedata                           (nios2cpu_data_master_writedata),                                        //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios2cpu_data_master_debugaccess),                                      //                          .debugaccess
		.i_address                             (nios2cpu_instruction_master_address),                                   //        instruction_master.address
		.i_read                                (nios2cpu_instruction_master_read),                                      //                          .read
		.i_readdata                            (nios2cpu_instruction_master_readdata),                                  //                          .readdata
		.i_waitrequest                         (nios2cpu_instruction_master_waitrequest),                               //                          .waitrequest
		.d_irq                                 (nios2cpu_d_irq_irq),                                                    //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2cpu_jtag_debug_module_reset_reset),                                //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_read),        //                          .read
		.jtag_debug_module_readdata            (nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_write),       //                          .write
		.jtag_debug_module_writedata           (nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                                       // custom_instruction_master.readra
	);

	DE0Qsys_sdram_ctrl sdram_ctrl (
		.clk            (syspll_c0_clk),                                              //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),                        // reset.reset_n
		.az_addr        (sdram_ctrl_s1_translator_avalon_anti_slave_0_address),       //    s1.address
		.az_be_n        (~sdram_ctrl_s1_translator_avalon_anti_slave_0_byteenable),   //      .byteenable_n
		.az_cs          (sdram_ctrl_s1_translator_avalon_anti_slave_0_chipselect),    //      .chipselect
		.az_data        (sdram_ctrl_s1_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.az_rd_n        (~sdram_ctrl_s1_translator_avalon_anti_slave_0_read),         //      .read_n
		.az_wr_n        (~sdram_ctrl_s1_translator_avalon_anti_slave_0_write),        //      .write_n
		.za_data        (sdram_ctrl_s1_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.za_valid       (sdram_ctrl_s1_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.za_waitrequest (sdram_ctrl_s1_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wires_addr),                                           //  wire.export
		.zs_ba          (sdram_wires_ba),                                             //      .export
		.zs_cas_n       (sdram_wires_cas_n),                                          //      .export
		.zs_cke         (sdram_wires_cke),                                            //      .export
		.zs_cs_n        (sdram_wires_cs_n),                                           //      .export
		.zs_dq          (sdram_wires_dq),                                             //      .export
		.zs_dqm         (sdram_wires_dqm),                                            //      .export
		.zs_ras_n       (sdram_wires_ras_n),                                          //      .export
		.zs_we_n        (sdram_wires_we_n)                                            //      .export
	);

	DE0Qsys_dma dma (
		.clk                (syspll_c0_clk),                                                    //                clk.clk
		.system_reset_n     (~rst_controller_001_reset_out_reset),                              //              reset.reset_n
		.dma_ctl_address    (dma_control_port_slave_translator_avalon_anti_slave_0_address),    // control_port_slave.address
		.dma_ctl_chipselect (dma_control_port_slave_translator_avalon_anti_slave_0_chipselect), //                   .chipselect
		.dma_ctl_readdata   (dma_control_port_slave_translator_avalon_anti_slave_0_readdata),   //                   .readdata
		.dma_ctl_write_n    (~dma_control_port_slave_translator_avalon_anti_slave_0_write),     //                   .write_n
		.dma_ctl_writedata  (dma_control_port_slave_translator_avalon_anti_slave_0_writedata),  //                   .writedata
		.dma_ctl_irq        (irq_mapper_receiver0_irq),                                         //                irq.irq
		.read_address       (dma_read_master_address),                                          //        read_master.address
		.read_chipselect    (dma_read_master_chipselect),                                       //                   .chipselect
		.read_read_n        (dma_read_master_read),                                             //                   .read_n
		.read_readdata      (dma_read_master_readdata),                                         //                   .readdata
		.read_readdatavalid (dma_read_master_readdatavalid),                                    //                   .readdatavalid
		.read_waitrequest   (dma_read_master_waitrequest),                                      //                   .waitrequest
		.read_burstcount    (dma_read_master_burstcount),                                       //                   .burstcount
		.write_address      (dma_write_master_address),                                         //       write_master.address
		.write_chipselect   (dma_write_master_chipselect),                                      //                   .chipselect
		.write_waitrequest  (dma_write_master_waitrequest),                                     //                   .waitrequest
		.write_write_n      (dma_write_master_write),                                           //                   .write_n
		.write_writedata    (dma_write_master_writedata),                                       //                   .writedata
		.write_byteenable   (dma_write_master_byteenable),                                      //                   .byteenable
		.write_burstcount   (dma_write_master_burstcount)                                       //                   .burstcount
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (10),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) apb (
		.clk              (syspll_c0_clk),                                       //   clk.clk
		.reset            (rst_controller_001_reset_out_reset),                  // reset.reset
		.s0_waitrequest   (apb_s0_translator_avalon_anti_slave_0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (apb_s0_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.s0_readdatavalid (apb_s0_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (apb_s0_translator_avalon_anti_slave_0_burstcount),    //      .burstcount
		.s0_writedata     (apb_s0_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.s0_address       (apb_s0_translator_avalon_anti_slave_0_address),       //      .address
		.s0_write         (apb_s0_translator_avalon_anti_slave_0_write),         //      .write
		.s0_read          (apb_s0_translator_avalon_anti_slave_0_read),          //      .read
		.s0_byteenable    (apb_s0_translator_avalon_anti_slave_0_byteenable),    //      .byteenable
		.s0_debugaccess   (apb_s0_translator_avalon_anti_slave_0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (apb_m0_waitrequest),                                  //    m0.waitrequest
		.m0_readdata      (apb_m0_readdata),                                     //      .readdata
		.m0_readdatavalid (apb_m0_readdatavalid),                                //      .readdatavalid
		.m0_burstcount    (apb_m0_burstcount),                                   //      .burstcount
		.m0_writedata     (apb_m0_writedata),                                    //      .writedata
		.m0_address       (apb_m0_address),                                      //      .address
		.m0_write         (apb_m0_write),                                        //      .write
		.m0_read          (apb_m0_read),                                         //      .read
		.m0_byteenable    (apb_m0_byteenable),                                   //      .byteenable
		.m0_debugaccess   (apb_m0_debugaccess)                                   //      .debugaccess
	);

	DE0Qsys_jtag_uart jtag_uart (
		.clk            (syspll_c0_clk),                                                          //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                                    //             reset.reset_n
		.av_chipselect  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                                //               irq.irq
	);

	DE0Qsys_timer timer (
		.clk        (syspll_c0_clk),                                      //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                // reset.reset_n
		.address    (timer_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                            //   irq.irq
	);

	DE0Qsys_uart0 uart0 (
		.clk           (syspll_c0_clk),                                         //                 clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),                   //               reset.reset_n
		.address       (uart0_s1_translator_avalon_anti_slave_0_address),       //                  s1.address
		.begintransfer (uart0_s1_translator_avalon_anti_slave_0_begintransfer), //                    .begintransfer
		.chipselect    (uart0_s1_translator_avalon_anti_slave_0_chipselect),    //                    .chipselect
		.read_n        (~uart0_s1_translator_avalon_anti_slave_0_read),         //                    .read_n
		.write_n       (~uart0_s1_translator_avalon_anti_slave_0_write),        //                    .write_n
		.writedata     (uart0_s1_translator_avalon_anti_slave_0_writedata),     //                    .writedata
		.readdata      (uart0_s1_translator_avalon_anti_slave_0_readdata),      //                    .readdata
		.dataavailable (),                                                      //                    .dataavailable
		.readyfordata  (),                                                      //                    .readyfordata
		.rxd           (uart0_rxd),                                             // external_connection.export
		.txd           (uart0_txd),                                             //                    .export
		.irq           (irq_mapper_receiver3_irq)                               //                 irq.irq
	);

	DE0Qsys_led led (
		.clk        (syspll_c0_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),              //               reset.reset_n
		.address    (led_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~led_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (led_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (led_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (led_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (led_export)                                        // external_connection.export
	);

	DE0Qsys_sw sw (
		.clk      (syspll_c0_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),           //               reset.reset_n
		.address  (sw_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (sw_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (sw_export)                                      // external_connection.export
	);

	DE0Qsys_button1 button1 (
		.clk        (syspll_c0_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                  //               reset.reset_n
		.address    (button1_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~button1_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (button1_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (button1_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (button1_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (button1_export),                                       // external_connection.export
		.irq        (irq_mapper_receiver4_irq)                              //                 irq.irq
	);

	DE0Qsys_button2 button2 (
		.clk      (syspll_c0_clk),                                      //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                //               reset.reset_n
		.address  (button2_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (button2_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (button2_export)                                      // external_connection.export
	);

	DE0Qsys_hex0 hex0 (
		.clk        (syspll_c0_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),               //               reset.reset_n
		.address    (hex0_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~hex0_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (hex0_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (hex0_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (hex0_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (hex0_export)                                        // external_connection.export
	);

	DE0Qsys_hex0 hex1 (
		.clk        (syspll_c0_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),               //               reset.reset_n
		.address    (hex1_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~hex1_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (hex1_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (hex1_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (hex1_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (hex1_export)                                        // external_connection.export
	);

	DE0Qsys_hex0 hex2 (
		.clk        (syspll_c0_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),               //               reset.reset_n
		.address    (hex2_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~hex2_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (hex2_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (hex2_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (hex2_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (hex2_export)                                        // external_connection.export
	);

	DE0Qsys_hex0 hex3 (
		.clk        (syspll_c0_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),               //               reset.reset_n
		.address    (hex3_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~hex3_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (hex3_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (hex3_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (hex3_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (hex3_export)                                        // external_connection.export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (26),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (26),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2cpu_instruction_master_translator (
		.clk                      (syspll_c0_clk),                                                                  //                       clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                             //                     reset.reset
		.uav_address              (nios2cpu_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (nios2cpu_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (nios2cpu_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (nios2cpu_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (nios2cpu_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (nios2cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (nios2cpu_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (nios2cpu_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (nios2cpu_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (nios2cpu_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (nios2cpu_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (nios2cpu_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (nios2cpu_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read                  (nios2cpu_instruction_master_read),                                               //                          .read
		.av_readdata              (nios2cpu_instruction_master_readdata),                                           //                          .readdata
		.av_burstcount            (1'b1),                                                                           //               (terminated)
		.av_byteenable            (4'b1111),                                                                        //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                           //               (terminated)
		.av_begintransfer         (1'b0),                                                                           //               (terminated)
		.av_chipselect            (1'b0),                                                                           //               (terminated)
		.av_readdatavalid         (),                                                                               //               (terminated)
		.av_write                 (1'b0),                                                                           //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                                           //               (terminated)
		.av_lock                  (1'b0),                                                                           //               (terminated)
		.av_debugaccess           (1'b0),                                                                           //               (terminated)
		.uav_clken                (),                                                                               //               (terminated)
		.av_clken                 (1'b1),                                                                           //               (terminated)
		.uav_response             (2'b00),                                                                          //               (terminated)
		.av_response              (),                                                                               //               (terminated)
		.uav_writeresponserequest (),                                                                               //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                           //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                           //               (terminated)
		.av_writeresponsevalid    ()                                                                                //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (26),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (8),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (26),
		.UAV_BURSTCOUNT_W            (10),
		.USE_READ                    (0),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (1),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (1),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) dma_write_master_translator (
		.clk                      (syspll_c0_clk),                                                       //                       clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                  //                     reset.reset
		.uav_address              (dma_write_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (dma_write_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (dma_write_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (dma_write_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (dma_write_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (dma_write_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (dma_write_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (dma_write_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (dma_write_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (dma_write_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (dma_write_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (dma_write_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (dma_write_master_waitrequest),                                        //                          .waitrequest
		.av_burstcount            (dma_write_master_burstcount),                                         //                          .burstcount
		.av_byteenable            (dma_write_master_byteenable),                                         //                          .byteenable
		.av_chipselect            (dma_write_master_chipselect),                                         //                          .chipselect
		.av_write                 (~dma_write_master_write),                                             //                          .write
		.av_writedata             (dma_write_master_writedata),                                          //                          .writedata
		.av_beginbursttransfer    (1'b0),                                                                //               (terminated)
		.av_begintransfer         (1'b0),                                                                //               (terminated)
		.av_read                  (1'b0),                                                                //               (terminated)
		.av_readdata              (),                                                                    //               (terminated)
		.av_readdatavalid         (),                                                                    //               (terminated)
		.av_lock                  (1'b0),                                                                //               (terminated)
		.av_debugaccess           (1'b0),                                                                //               (terminated)
		.uav_clken                (),                                                                    //               (terminated)
		.av_clken                 (1'b1),                                                                //               (terminated)
		.uav_response             (2'b00),                                                               //               (terminated)
		.av_response              (),                                                                    //               (terminated)
		.uav_writeresponserequest (),                                                                    //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                //               (terminated)
		.av_writeresponsevalid    ()                                                                     //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (26),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (26),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (1)
	) nios2cpu_data_master_translator (
		.clk                      (syspll_c0_clk),                                                           //                       clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                      //                     reset.reset
		.uav_address              (nios2cpu_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (nios2cpu_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (nios2cpu_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (nios2cpu_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (nios2cpu_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (nios2cpu_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (nios2cpu_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (nios2cpu_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (nios2cpu_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (nios2cpu_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (nios2cpu_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (nios2cpu_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (nios2cpu_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (nios2cpu_data_master_byteenable),                                         //                          .byteenable
		.av_read                  (nios2cpu_data_master_read),                                               //                          .read
		.av_readdata              (nios2cpu_data_master_readdata),                                           //                          .readdata
		.av_write                 (nios2cpu_data_master_write),                                              //                          .write
		.av_writedata             (nios2cpu_data_master_writedata),                                          //                          .writedata
		.av_debugaccess           (nios2cpu_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount            (1'b1),                                                                    //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                    //               (terminated)
		.av_begintransfer         (1'b0),                                                                    //               (terminated)
		.av_chipselect            (1'b0),                                                                    //               (terminated)
		.av_readdatavalid         (),                                                                        //               (terminated)
		.av_lock                  (1'b0),                                                                    //               (terminated)
		.uav_clken                (),                                                                        //               (terminated)
		.av_clken                 (1'b1),                                                                    //               (terminated)
		.uav_response             (2'b00),                                                                   //               (terminated)
		.av_response              (),                                                                        //               (terminated)
		.uav_writeresponserequest (),                                                                        //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                    //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                    //               (terminated)
		.av_writeresponsevalid    ()                                                                         //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (26),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (8),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (26),
		.UAV_BURSTCOUNT_W            (10),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (1),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (1),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) dma_read_master_translator (
		.clk                      (syspll_c0_clk),                                                      //                       clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                 //                     reset.reset
		.uav_address              (dma_read_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (dma_read_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (dma_read_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (dma_read_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (dma_read_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (dma_read_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (dma_read_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (dma_read_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (dma_read_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (dma_read_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (dma_read_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (dma_read_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (dma_read_master_waitrequest),                                        //                          .waitrequest
		.av_burstcount            (dma_read_master_burstcount),                                         //                          .burstcount
		.av_chipselect            (dma_read_master_chipselect),                                         //                          .chipselect
		.av_read                  (~dma_read_master_read),                                              //                          .read
		.av_readdata              (dma_read_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (dma_read_master_readdatavalid),                                      //                          .readdatavalid
		.av_byteenable            (4'b1111),                                                            //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                               //               (terminated)
		.av_begintransfer         (1'b0),                                                               //               (terminated)
		.av_write                 (1'b0),                                                               //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                               //               (terminated)
		.av_lock                  (1'b0),                                                               //               (terminated)
		.av_debugaccess           (1'b0),                                                               //               (terminated)
		.uav_clken                (),                                                                   //               (terminated)
		.av_clken                 (1'b1),                                                               //               (terminated)
		.uav_response             (2'b00),                                                              //               (terminated)
		.av_response              (),                                                                   //               (terminated)
		.uav_writeresponserequest (),                                                                   //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                               //               (terminated)
		.av_writeresponserequest  (1'b0),                                                               //               (terminated)
		.av_writeresponsevalid    ()                                                                    //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) nios2cpu_jtag_debug_module_translator (
		.clk                      (syspll_c0_clk),                                                                         //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                                    //                    reset.reset
		.uav_address              (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess           (nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                                      //              (terminated)
		.av_burstcount            (),                                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                                      //              (terminated)
		.av_lock                  (),                                                                                      //              (terminated)
		.av_chipselect            (),                                                                                      //              (terminated)
		.av_clken                 (),                                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                                  //              (terminated)
		.av_outputenable          (),                                                                                      //              (terminated)
		.uav_response             (),                                                                                      //              (terminated)
		.av_response              (2'b00),                                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (22),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sdram_ctrl_s1_translator (
		.clk                      (syspll_c0_clk),                                                            //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sdram_ctrl_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (sdram_ctrl_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (sdram_ctrl_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (sdram_ctrl_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (sdram_ctrl_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (sdram_ctrl_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (sdram_ctrl_s1_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (sdram_ctrl_s1_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (sdram_ctrl_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (26),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) dma_control_port_slave_translator (
		.clk                      (syspll_c0_clk),                                                                     //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                                //                    reset.reset
		.uav_address              (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (dma_control_port_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (dma_control_port_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (dma_control_port_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (dma_control_port_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (dma_control_port_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                                  //              (terminated)
		.av_begintransfer         (),                                                                                  //              (terminated)
		.av_beginbursttransfer    (),                                                                                  //              (terminated)
		.av_burstcount            (),                                                                                  //              (terminated)
		.av_byteenable            (),                                                                                  //              (terminated)
		.av_readdatavalid         (1'b0),                                                                              //              (terminated)
		.av_waitrequest           (1'b0),                                                                              //              (terminated)
		.av_writebyteenable       (),                                                                                  //              (terminated)
		.av_lock                  (),                                                                                  //              (terminated)
		.av_clken                 (),                                                                                  //              (terminated)
		.uav_clken                (1'b0),                                                                              //              (terminated)
		.av_debugaccess           (),                                                                                  //              (terminated)
		.av_outputenable          (),                                                                                  //              (terminated)
		.uav_response             (),                                                                                  //              (terminated)
		.av_response              (2'b00),                                                                             //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                              //              (terminated)
		.uav_writeresponsevalid   (),                                                                                  //              (terminated)
		.av_writeresponserequest  (),                                                                                  //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (10),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) apb_s0_translator (
		.clk                      (syspll_c0_clk),                                                     //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                //                    reset.reset
		.uav_address              (apb_s0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (apb_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (apb_s0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (apb_s0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (apb_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (apb_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (apb_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (apb_s0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (apb_s0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (apb_s0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (apb_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (apb_s0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (apb_s0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (apb_s0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (apb_s0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (apb_s0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount            (apb_s0_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable            (apb_s0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (apb_s0_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (apb_s0_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess           (apb_s0_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                  //              (terminated)
		.av_beginbursttransfer    (),                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                  //              (terminated)
		.av_lock                  (),                                                                  //              (terminated)
		.av_chipselect            (),                                                                  //              (terminated)
		.av_clken                 (),                                                                  //              (terminated)
		.uav_clken                (1'b0),                                                              //              (terminated)
		.av_outputenable          (),                                                                  //              (terminated)
		.uav_response             (),                                                                  //              (terminated)
		.av_response              (2'b00),                                                             //              (terminated)
		.uav_writeresponserequest (1'b0),                                                              //              (terminated)
		.uav_writeresponsevalid   (),                                                                  //              (terminated)
		.av_writeresponserequest  (),                                                                  //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) syspll_pll_slave_translator (
		.clk                      (clk_50m_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                              //                    reset.reset
		.uav_address              (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (syspll_pll_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (syspll_pll_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (syspll_pll_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (syspll_pll_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (syspll_pll_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (),                                                                            //              (terminated)
		.av_beginbursttransfer    (),                                                                            //              (terminated)
		.av_burstcount            (),                                                                            //              (terminated)
		.av_byteenable            (),                                                                            //              (terminated)
		.av_readdatavalid         (1'b0),                                                                        //              (terminated)
		.av_waitrequest           (1'b0),                                                                        //              (terminated)
		.av_writebyteenable       (),                                                                            //              (terminated)
		.av_lock                  (),                                                                            //              (terminated)
		.av_chipselect            (),                                                                            //              (terminated)
		.av_clken                 (),                                                                            //              (terminated)
		.uav_clken                (1'b0),                                                                        //              (terminated)
		.av_debugaccess           (),                                                                            //              (terminated)
		.av_outputenable          (),                                                                            //              (terminated)
		.uav_response             (),                                                                            //              (terminated)
		.av_response              (2'b00),                                                                       //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                        //              (terminated)
		.uav_writeresponsevalid   (),                                                                            //              (terminated)
		.av_writeresponserequest  (),                                                                            //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                         //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (10),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (10),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) apb_m0_translator (
		.clk                      (syspll_c0_clk),                                             //                       clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                        //                     reset.reset
		.uav_address              (apb_m0_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (apb_m0_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (apb_m0_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (apb_m0_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (apb_m0_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (apb_m0_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (apb_m0_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (apb_m0_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (apb_m0_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (apb_m0_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (apb_m0_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (apb_m0_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (apb_m0_waitrequest),                                        //                          .waitrequest
		.av_burstcount            (apb_m0_burstcount),                                         //                          .burstcount
		.av_byteenable            (apb_m0_byteenable),                                         //                          .byteenable
		.av_read                  (apb_m0_read),                                               //                          .read
		.av_readdata              (apb_m0_readdata),                                           //                          .readdata
		.av_readdatavalid         (apb_m0_readdatavalid),                                      //                          .readdatavalid
		.av_write                 (apb_m0_write),                                              //                          .write
		.av_writedata             (apb_m0_writedata),                                          //                          .writedata
		.av_debugaccess           (apb_m0_debugaccess),                                        //                          .debugaccess
		.av_beginbursttransfer    (1'b0),                                                      //               (terminated)
		.av_begintransfer         (1'b0),                                                      //               (terminated)
		.av_chipselect            (1'b0),                                                      //               (terminated)
		.av_lock                  (1'b0),                                                      //               (terminated)
		.uav_clken                (),                                                          //               (terminated)
		.av_clken                 (1'b1),                                                      //               (terminated)
		.uav_response             (2'b00),                                                     //               (terminated)
		.av_response              (),                                                          //               (terminated)
		.uav_writeresponserequest (),                                                          //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                      //               (terminated)
		.av_writeresponserequest  (1'b0),                                                      //               (terminated)
		.av_writeresponsevalid    ()                                                           //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_avalon_jtag_slave_translator (
		.clk                      (syspll_c0_clk),                                                                          //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                                     //                    reset.reset
		.uav_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                                       //              (terminated)
		.av_burstcount            (),                                                                                       //              (terminated)
		.av_byteenable            (),                                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                                       //              (terminated)
		.av_lock                  (),                                                                                       //              (terminated)
		.av_clken                 (),                                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                                   //              (terminated)
		.av_debugaccess           (),                                                                                       //              (terminated)
		.av_outputenable          (),                                                                                       //              (terminated)
		.uav_response             (),                                                                                       //              (terminated)
		.av_response              (2'b00),                                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_s1_translator (
		.clk                      (syspll_c0_clk),                                                       //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                  //                    reset.reset
		.uav_address              (timer_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (timer_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (timer_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (timer_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (timer_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (timer_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (timer_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (timer_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                    //              (terminated)
		.av_begintransfer         (),                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                    //              (terminated)
		.av_burstcount            (),                                                                    //              (terminated)
		.av_byteenable            (),                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                //              (terminated)
		.av_waitrequest           (1'b0),                                                                //              (terminated)
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) uart0_s1_translator (
		.clk                      (syspll_c0_clk),                                                       //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                  //                    reset.reset
		.uav_address              (uart0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (uart0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (uart0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (uart0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (uart0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (uart0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (uart0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (uart0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (uart0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (uart0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (uart0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (uart0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (uart0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (uart0_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (uart0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (uart0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (uart0_s1_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_chipselect            (uart0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_beginbursttransfer    (),                                                                    //              (terminated)
		.av_burstcount            (),                                                                    //              (terminated)
		.av_byteenable            (),                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                //              (terminated)
		.av_waitrequest           (1'b0),                                                                //              (terminated)
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sw_s1_translator (
		.clk                      (syspll_c0_clk),                                                    //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                               //                    reset.reset
		.uav_address              (sw_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sw_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sw_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sw_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sw_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sw_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sw_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sw_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sw_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sw_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sw_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sw_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (sw_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                 //              (terminated)
		.av_read                  (),                                                                 //              (terminated)
		.av_writedata             (),                                                                 //              (terminated)
		.av_begintransfer         (),                                                                 //              (terminated)
		.av_beginbursttransfer    (),                                                                 //              (terminated)
		.av_burstcount            (),                                                                 //              (terminated)
		.av_byteenable            (),                                                                 //              (terminated)
		.av_readdatavalid         (1'b0),                                                             //              (terminated)
		.av_waitrequest           (1'b0),                                                             //              (terminated)
		.av_writebyteenable       (),                                                                 //              (terminated)
		.av_lock                  (),                                                                 //              (terminated)
		.av_chipselect            (),                                                                 //              (terminated)
		.av_clken                 (),                                                                 //              (terminated)
		.uav_clken                (1'b0),                                                             //              (terminated)
		.av_debugaccess           (),                                                                 //              (terminated)
		.av_outputenable          (),                                                                 //              (terminated)
		.uav_response             (),                                                                 //              (terminated)
		.av_response              (2'b00),                                                            //              (terminated)
		.uav_writeresponserequest (1'b0),                                                             //              (terminated)
		.uav_writeresponsevalid   (),                                                                 //              (terminated)
		.av_writeresponserequest  (),                                                                 //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) led_s1_translator (
		.clk                      (syspll_c0_clk),                                                     //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                //                    reset.reset
		.uav_address              (led_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (led_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (led_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (led_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (led_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (led_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (led_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (led_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (led_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (led_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (led_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (led_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (led_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (led_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (led_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (led_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                  //              (terminated)
		.av_begintransfer         (),                                                                  //              (terminated)
		.av_beginbursttransfer    (),                                                                  //              (terminated)
		.av_burstcount            (),                                                                  //              (terminated)
		.av_byteenable            (),                                                                  //              (terminated)
		.av_readdatavalid         (1'b0),                                                              //              (terminated)
		.av_waitrequest           (1'b0),                                                              //              (terminated)
		.av_writebyteenable       (),                                                                  //              (terminated)
		.av_lock                  (),                                                                  //              (terminated)
		.av_clken                 (),                                                                  //              (terminated)
		.uav_clken                (1'b0),                                                              //              (terminated)
		.av_debugaccess           (),                                                                  //              (terminated)
		.av_outputenable          (),                                                                  //              (terminated)
		.uav_response             (),                                                                  //              (terminated)
		.av_response              (2'b00),                                                             //              (terminated)
		.uav_writeresponserequest (1'b0),                                                              //              (terminated)
		.uav_writeresponsevalid   (),                                                                  //              (terminated)
		.av_writeresponserequest  (),                                                                  //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) button1_s1_translator (
		.clk                      (syspll_c0_clk),                                                         //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                    //                    reset.reset
		.uav_address              (button1_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (button1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (button1_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (button1_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (button1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (button1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (button1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (button1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (button1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (button1_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (button1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (button1_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (button1_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (button1_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (button1_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (button1_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                      //              (terminated)
		.av_begintransfer         (),                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                      //              (terminated)
		.av_burstcount            (),                                                                      //              (terminated)
		.av_byteenable            (),                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                      //              (terminated)
		.av_lock                  (),                                                                      //              (terminated)
		.av_clken                 (),                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                  //              (terminated)
		.av_debugaccess           (),                                                                      //              (terminated)
		.av_outputenable          (),                                                                      //              (terminated)
		.uav_response             (),                                                                      //              (terminated)
		.av_response              (2'b00),                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) button2_s1_translator (
		.clk                      (syspll_c0_clk),                                                         //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                    //                    reset.reset
		.uav_address              (button2_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (button2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (button2_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (button2_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (button2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (button2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (button2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (button2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (button2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (button2_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (button2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (button2_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (button2_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                      //              (terminated)
		.av_read                  (),                                                                      //              (terminated)
		.av_writedata             (),                                                                      //              (terminated)
		.av_begintransfer         (),                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                      //              (terminated)
		.av_burstcount            (),                                                                      //              (terminated)
		.av_byteenable            (),                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                      //              (terminated)
		.av_lock                  (),                                                                      //              (terminated)
		.av_chipselect            (),                                                                      //              (terminated)
		.av_clken                 (),                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                  //              (terminated)
		.av_debugaccess           (),                                                                      //              (terminated)
		.av_outputenable          (),                                                                      //              (terminated)
		.uav_response             (),                                                                      //              (terminated)
		.av_response              (2'b00),                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) hex0_s1_translator (
		.clk                      (syspll_c0_clk),                                                      //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                 //                    reset.reset
		.uav_address              (hex0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (hex0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (hex0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (hex0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (hex0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (hex0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (hex0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (hex0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (hex0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (hex0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (hex0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (hex0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (hex0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (hex0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (hex0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (hex0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                   //              (terminated)
		.av_begintransfer         (),                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                   //              (terminated)
		.av_burstcount            (),                                                                   //              (terminated)
		.av_byteenable            (),                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                               //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) hex1_s1_translator (
		.clk                      (syspll_c0_clk),                                                      //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                 //                    reset.reset
		.uav_address              (hex1_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (hex1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (hex1_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (hex1_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (hex1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (hex1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (hex1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (hex1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (hex1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (hex1_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (hex1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (hex1_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (hex1_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (hex1_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (hex1_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (hex1_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                   //              (terminated)
		.av_begintransfer         (),                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                   //              (terminated)
		.av_burstcount            (),                                                                   //              (terminated)
		.av_byteenable            (),                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                               //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) hex2_s1_translator (
		.clk                      (syspll_c0_clk),                                                      //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                 //                    reset.reset
		.uav_address              (hex2_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (hex2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (hex2_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (hex2_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (hex2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (hex2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (hex2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (hex2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (hex2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (hex2_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (hex2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (hex2_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (hex2_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (hex2_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (hex2_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (hex2_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                   //              (terminated)
		.av_begintransfer         (),                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                   //              (terminated)
		.av_burstcount            (),                                                                   //              (terminated)
		.av_byteenable            (),                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                               //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) hex3_s1_translator (
		.clk                      (syspll_c0_clk),                                                      //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                 //                    reset.reset
		.uav_address              (hex3_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (hex3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (hex3_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (hex3_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (hex3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (hex3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (hex3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (hex3_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (hex3_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (hex3_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (hex3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (hex3_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (hex3_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (hex3_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (hex3_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (hex3_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                   //              (terminated)
		.av_begintransfer         (),                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                   //              (terminated)
		.av_burstcount            (),                                                                   //              (terminated)
		.av_byteenable            (),                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                               //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (99),
		.PKT_PROTECTION_L          (97),
		.PKT_BEGIN_BURST           (88),
		.PKT_BURSTWRAP_H           (80),
		.PKT_BURSTWRAP_L           (78),
		.PKT_BURST_SIZE_H          (83),
		.PKT_BURST_SIZE_L          (81),
		.PKT_BURST_TYPE_H          (85),
		.PKT_BURST_TYPE_L          (84),
		.PKT_BYTE_CNT_H            (77),
		.PKT_BYTE_CNT_L            (68),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_TRANS_EXCLUSIVE       (67),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (90),
		.PKT_DEST_ID_H             (95),
		.PKT_DEST_ID_L             (93),
		.PKT_THREAD_ID_H           (96),
		.PKT_THREAD_ID_L           (96),
		.PKT_CACHE_H               (103),
		.PKT_CACHE_L               (100),
		.PKT_DATA_SIDEBAND_H       (87),
		.PKT_DATA_SIDEBAND_L       (87),
		.PKT_QOS_H                 (89),
		.PKT_QOS_L                 (89),
		.PKT_ADDR_SIDEBAND_H       (86),
		.PKT_ADDR_SIDEBAND_L       (86),
		.PKT_RESPONSE_STATUS_H     (105),
		.PKT_RESPONSE_STATUS_L     (104),
		.ST_DATA_W                 (106),
		.ST_CHANNEL_W              (5),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (3),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2cpu_instruction_master_translator_avalon_universal_master_0_agent (
		.clk                     (syspll_c0_clk),                                                                           //       clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                      // clk_reset.reset
		.av_address              (nios2cpu_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (nios2cpu_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (nios2cpu_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (nios2cpu_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (nios2cpu_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (nios2cpu_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (nios2cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (nios2cpu_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (nios2cpu_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (nios2cpu_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (nios2cpu_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (nios2cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (nios2cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (nios2cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (nios2cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (nios2cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_src_valid),                                                                  //        rp.valid
		.rp_data                 (rsp_xbar_mux_src_data),                                                                   //          .data
		.rp_channel              (rsp_xbar_mux_src_channel),                                                                //          .channel
		.rp_startofpacket        (rsp_xbar_mux_src_startofpacket),                                                          //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_src_endofpacket),                                                            //          .endofpacket
		.rp_ready                (rsp_xbar_mux_src_ready),                                                                  //          .ready
		.av_response             (),                                                                                        // (terminated)
		.av_writeresponserequest (1'b0),                                                                                    // (terminated)
		.av_writeresponsevalid   ()                                                                                         // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (99),
		.PKT_PROTECTION_L          (97),
		.PKT_BEGIN_BURST           (88),
		.PKT_BURSTWRAP_H           (80),
		.PKT_BURSTWRAP_L           (78),
		.PKT_BURST_SIZE_H          (83),
		.PKT_BURST_SIZE_L          (81),
		.PKT_BURST_TYPE_H          (85),
		.PKT_BURST_TYPE_L          (84),
		.PKT_BYTE_CNT_H            (77),
		.PKT_BYTE_CNT_L            (68),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_TRANS_EXCLUSIVE       (67),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (90),
		.PKT_DEST_ID_H             (95),
		.PKT_DEST_ID_L             (93),
		.PKT_THREAD_ID_H           (96),
		.PKT_THREAD_ID_L           (96),
		.PKT_CACHE_H               (103),
		.PKT_CACHE_L               (100),
		.PKT_DATA_SIDEBAND_H       (87),
		.PKT_DATA_SIDEBAND_L       (87),
		.PKT_QOS_H                 (89),
		.PKT_QOS_L                 (89),
		.PKT_ADDR_SIDEBAND_H       (86),
		.PKT_ADDR_SIDEBAND_L       (86),
		.PKT_RESPONSE_STATUS_H     (105),
		.PKT_RESPONSE_STATUS_L     (104),
		.ST_DATA_W                 (106),
		.ST_CHANNEL_W              (5),
		.AV_BURSTCOUNT_W           (10),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) dma_write_master_translator_avalon_universal_master_0_agent (
		.clk                     (syspll_c0_clk),                                                                //       clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.av_address              (dma_write_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (dma_write_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (dma_write_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (dma_write_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (dma_write_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (dma_write_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (dma_write_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (dma_write_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (dma_write_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (dma_write_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (dma_write_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (dma_write_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (dma_write_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (dma_write_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (dma_write_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (dma_write_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_001_src_valid),                                                   //        rp.valid
		.rp_data                 (rsp_xbar_mux_001_src_data),                                                    //          .data
		.rp_channel              (rsp_xbar_mux_001_src_channel),                                                 //          .channel
		.rp_startofpacket        (rsp_xbar_mux_001_src_startofpacket),                                           //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_001_src_endofpacket),                                             //          .endofpacket
		.rp_ready                (rsp_xbar_mux_001_src_ready),                                                   //          .ready
		.av_response             (),                                                                             // (terminated)
		.av_writeresponserequest (1'b0),                                                                         // (terminated)
		.av_writeresponsevalid   ()                                                                              // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (99),
		.PKT_PROTECTION_L          (97),
		.PKT_BEGIN_BURST           (88),
		.PKT_BURSTWRAP_H           (80),
		.PKT_BURSTWRAP_L           (78),
		.PKT_BURST_SIZE_H          (83),
		.PKT_BURST_SIZE_L          (81),
		.PKT_BURST_TYPE_H          (85),
		.PKT_BURST_TYPE_L          (84),
		.PKT_BYTE_CNT_H            (77),
		.PKT_BYTE_CNT_L            (68),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_TRANS_EXCLUSIVE       (67),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (90),
		.PKT_DEST_ID_H             (95),
		.PKT_DEST_ID_L             (93),
		.PKT_THREAD_ID_H           (96),
		.PKT_THREAD_ID_L           (96),
		.PKT_CACHE_H               (103),
		.PKT_CACHE_L               (100),
		.PKT_DATA_SIDEBAND_H       (87),
		.PKT_DATA_SIDEBAND_L       (87),
		.PKT_QOS_H                 (89),
		.PKT_QOS_L                 (89),
		.PKT_ADDR_SIDEBAND_H       (86),
		.PKT_ADDR_SIDEBAND_L       (86),
		.PKT_RESPONSE_STATUS_H     (105),
		.PKT_RESPONSE_STATUS_L     (104),
		.ST_DATA_W                 (106),
		.ST_CHANNEL_W              (5),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (2),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2cpu_data_master_translator_avalon_universal_master_0_agent (
		.clk                     (syspll_c0_clk),                                                                    //       clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                               // clk_reset.reset
		.av_address              (nios2cpu_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (nios2cpu_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (nios2cpu_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (nios2cpu_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (nios2cpu_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (nios2cpu_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (nios2cpu_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (nios2cpu_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (nios2cpu_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (nios2cpu_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (nios2cpu_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (nios2cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (nios2cpu_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (nios2cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (nios2cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (nios2cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_002_src_valid),                                                       //        rp.valid
		.rp_data                 (rsp_xbar_mux_002_src_data),                                                        //          .data
		.rp_channel              (rsp_xbar_mux_002_src_channel),                                                     //          .channel
		.rp_startofpacket        (rsp_xbar_mux_002_src_startofpacket),                                               //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_002_src_endofpacket),                                                 //          .endofpacket
		.rp_ready                (rsp_xbar_mux_002_src_ready),                                                       //          .ready
		.av_response             (),                                                                                 // (terminated)
		.av_writeresponserequest (1'b0),                                                                             // (terminated)
		.av_writeresponsevalid   ()                                                                                  // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (99),
		.PKT_PROTECTION_L          (97),
		.PKT_BEGIN_BURST           (88),
		.PKT_BURSTWRAP_H           (80),
		.PKT_BURSTWRAP_L           (78),
		.PKT_BURST_SIZE_H          (83),
		.PKT_BURST_SIZE_L          (81),
		.PKT_BURST_TYPE_H          (85),
		.PKT_BURST_TYPE_L          (84),
		.PKT_BYTE_CNT_H            (77),
		.PKT_BYTE_CNT_L            (68),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_TRANS_EXCLUSIVE       (67),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (90),
		.PKT_DEST_ID_H             (95),
		.PKT_DEST_ID_L             (93),
		.PKT_THREAD_ID_H           (96),
		.PKT_THREAD_ID_L           (96),
		.PKT_CACHE_H               (103),
		.PKT_CACHE_L               (100),
		.PKT_DATA_SIDEBAND_H       (87),
		.PKT_DATA_SIDEBAND_L       (87),
		.PKT_QOS_H                 (89),
		.PKT_QOS_L                 (89),
		.PKT_ADDR_SIDEBAND_H       (86),
		.PKT_ADDR_SIDEBAND_L       (86),
		.PKT_RESPONSE_STATUS_H     (105),
		.PKT_RESPONSE_STATUS_L     (104),
		.ST_DATA_W                 (106),
		.ST_CHANNEL_W              (5),
		.AV_BURSTCOUNT_W           (10),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) dma_read_master_translator_avalon_universal_master_0_agent (
		.clk                     (syspll_c0_clk),                                                               //       clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.av_address              (dma_read_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (dma_read_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (dma_read_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (dma_read_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (dma_read_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (dma_read_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (dma_read_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (dma_read_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (dma_read_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (dma_read_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (dma_read_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (dma_read_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (dma_read_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (dma_read_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (dma_read_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (dma_read_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (limiter_rsp_src_valid),                                                       //        rp.valid
		.rp_data                 (limiter_rsp_src_data),                                                        //          .data
		.rp_channel              (limiter_rsp_src_channel),                                                     //          .channel
		.rp_startofpacket        (limiter_rsp_src_startofpacket),                                               //          .startofpacket
		.rp_endofpacket          (limiter_rsp_src_endofpacket),                                                 //          .endofpacket
		.rp_ready                (limiter_rsp_src_ready),                                                       //          .ready
		.av_response             (),                                                                            // (terminated)
		.av_writeresponserequest (1'b0),                                                                        // (terminated)
		.av_writeresponsevalid   ()                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (88),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (90),
		.PKT_DEST_ID_H             (95),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (80),
		.PKT_BURSTWRAP_L           (78),
		.PKT_BYTE_CNT_H            (77),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (99),
		.PKT_PROTECTION_L          (97),
		.PKT_RESPONSE_STATUS_H     (105),
		.PKT_RESPONSE_STATUS_L     (104),
		.PKT_BURST_SIZE_H          (83),
		.PKT_BURST_SIZE_L          (81),
		.ST_CHANNEL_W              (5),
		.ST_DATA_W                 (106),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (syspll_c0_clk),                                                                                   //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                              //       clk_reset.reset
		.m0_address              (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                          //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                          //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                           //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                                  //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                                    //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                        //                .channel
		.rf_sink_ready           (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (107),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (syspll_c0_clk),                                                                                   //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                              // clk_reset.reset
		.in_data           (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                           // (terminated)
		.csr_read          (1'b0),                                                                                            // (terminated)
		.csr_write         (1'b0),                                                                                            // (terminated)
		.csr_readdata      (),                                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                            // (terminated)
		.almost_full_data  (),                                                                                                // (terminated)
		.almost_empty_data (),                                                                                                // (terminated)
		.in_empty          (1'b0),                                                                                            // (terminated)
		.out_empty         (),                                                                                                // (terminated)
		.in_error          (1'b0),                                                                                            // (terminated)
		.out_error         (),                                                                                                // (terminated)
		.in_channel        (1'b0),                                                                                            // (terminated)
		.out_channel       ()                                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (70),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (43),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (44),
		.PKT_TRANS_POSTED          (45),
		.PKT_TRANS_WRITE           (46),
		.PKT_TRANS_READ            (47),
		.PKT_TRANS_LOCK            (48),
		.PKT_SRC_ID_H              (74),
		.PKT_SRC_ID_L              (72),
		.PKT_DEST_ID_H             (77),
		.PKT_DEST_ID_L             (75),
		.PKT_BURSTWRAP_H           (62),
		.PKT_BURSTWRAP_L           (60),
		.PKT_BYTE_CNT_H            (59),
		.PKT_BYTE_CNT_L            (50),
		.PKT_PROTECTION_H          (81),
		.PKT_PROTECTION_L          (79),
		.PKT_RESPONSE_STATUS_H     (87),
		.PKT_RESPONSE_STATUS_L     (86),
		.PKT_BURST_SIZE_H          (65),
		.PKT_BURST_SIZE_L          (63),
		.ST_CHANNEL_W              (5),
		.ST_DATA_W                 (88),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sdram_ctrl_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (syspll_c0_clk),                                                                      //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                        //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                        //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                         //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                                  //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                      //                .channel
		.rf_sink_ready           (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (89),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (syspll_c0_clk),                                                                      //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (18),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (syspll_c0_clk),                                                                //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.in_data           (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_startofpacket  (1'b0),                                                                         // (terminated)
		.in_endofpacket    (1'b0),                                                                         // (terminated)
		.out_startofpacket (),                                                                             // (terminated)
		.out_endofpacket   (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (88),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (90),
		.PKT_DEST_ID_H             (95),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (80),
		.PKT_BURSTWRAP_L           (78),
		.PKT_BYTE_CNT_H            (77),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (99),
		.PKT_PROTECTION_L          (97),
		.PKT_RESPONSE_STATUS_H     (105),
		.PKT_RESPONSE_STATUS_L     (104),
		.PKT_BURST_SIZE_H          (83),
		.PKT_BURST_SIZE_L          (81),
		.ST_CHANNEL_W              (5),
		.ST_DATA_W                 (106),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) dma_control_port_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (syspll_c0_clk),                                                                               //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                          //       clk_reset.reset
		.m0_address              (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_002_src_ready),                                                                  //              cp.ready
		.cp_valid                (cmd_xbar_mux_002_src_valid),                                                                  //                .valid
		.cp_data                 (cmd_xbar_mux_002_src_data),                                                                   //                .data
		.cp_startofpacket        (cmd_xbar_mux_002_src_startofpacket),                                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_002_src_endofpacket),                                                            //                .endofpacket
		.cp_channel              (cmd_xbar_mux_002_src_channel),                                                                //                .channel
		.rf_sink_ready           (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                       //     (terminated)
		.m0_writeresponserequest (),                                                                                            //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                         //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (107),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (syspll_c0_clk),                                                                               //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                          // clk_reset.reset
		.in_data           (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                        // (terminated)
		.csr_readdata      (),                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                        // (terminated)
		.almost_full_data  (),                                                                                            // (terminated)
		.almost_empty_data (),                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                        // (terminated)
		.out_empty         (),                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                        // (terminated)
		.out_error         (),                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                        // (terminated)
		.out_channel       ()                                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (88),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (90),
		.PKT_DEST_ID_H             (95),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (80),
		.PKT_BURSTWRAP_L           (78),
		.PKT_BYTE_CNT_H            (77),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (99),
		.PKT_PROTECTION_L          (97),
		.PKT_RESPONSE_STATUS_H     (105),
		.PKT_RESPONSE_STATUS_L     (104),
		.PKT_BURST_SIZE_H          (83),
		.PKT_BURST_SIZE_L          (81),
		.ST_CHANNEL_W              (5),
		.ST_DATA_W                 (106),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) apb_s0_translator_avalon_universal_slave_0_agent (
		.clk                     (syspll_c0_clk),                                                               //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                          //       clk_reset.reset
		.m0_address              (apb_s0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (apb_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (apb_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (apb_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (apb_s0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (apb_s0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (apb_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (apb_s0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (apb_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (apb_s0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (apb_s0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (apb_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (apb_s0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (apb_s0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (apb_s0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (apb_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_001_source0_ready),                                             //              cp.ready
		.cp_valid                (burst_adapter_001_source0_valid),                                             //                .valid
		.cp_data                 (burst_adapter_001_source0_data),                                              //                .data
		.cp_startofpacket        (burst_adapter_001_source0_startofpacket),                                     //                .startofpacket
		.cp_endofpacket          (burst_adapter_001_source0_endofpacket),                                       //                .endofpacket
		.cp_channel              (burst_adapter_001_source0_channel),                                           //                .channel
		.rf_sink_ready           (apb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (apb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (apb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (apb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (apb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (apb_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (apb_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (apb_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (apb_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (apb_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (apb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (apb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (apb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (apb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (apb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (apb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                       //     (terminated)
		.m0_writeresponserequest (),                                                                            //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                         //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (107),
		.FIFO_DEPTH          (5),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) apb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (syspll_c0_clk),                                                               //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.in_data           (apb_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (apb_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (apb_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (apb_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (apb_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (apb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (apb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (apb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (apb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (apb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                       // (terminated)
		.csr_read          (1'b0),                                                                        // (terminated)
		.csr_write         (1'b0),                                                                        // (terminated)
		.csr_readdata      (),                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                        // (terminated)
		.almost_full_data  (),                                                                            // (terminated)
		.almost_empty_data (),                                                                            // (terminated)
		.in_empty          (1'b0),                                                                        // (terminated)
		.out_empty         (),                                                                            // (terminated)
		.in_error          (1'b0),                                                                        // (terminated)
		.out_error         (),                                                                            // (terminated)
		.in_channel        (1'b0),                                                                        // (terminated)
		.out_channel       ()                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (88),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (90),
		.PKT_DEST_ID_H             (95),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (80),
		.PKT_BURSTWRAP_L           (78),
		.PKT_BYTE_CNT_H            (77),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (99),
		.PKT_PROTECTION_L          (97),
		.PKT_RESPONSE_STATUS_H     (105),
		.PKT_RESPONSE_STATUS_L     (104),
		.PKT_BURST_SIZE_H          (83),
		.PKT_BURST_SIZE_L          (81),
		.ST_CHANNEL_W              (5),
		.ST_DATA_W                 (106),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) syspll_pll_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_50m_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_out_ready),                                                                     //              cp.ready
		.cp_valid                (crosser_out_valid),                                                                     //                .valid
		.cp_data                 (crosser_out_data),                                                                      //                .data
		.cp_startofpacket        (crosser_out_startofpacket),                                                             //                .startofpacket
		.cp_endofpacket          (crosser_out_endofpacket),                                                               //                .endofpacket
		.cp_channel              (crosser_out_channel),                                                                   //                .channel
		.rf_sink_ready           (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                 //     (terminated)
		.m0_writeresponserequest (),                                                                                      //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                   //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (107),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_50m_clk),                                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_50m_clk),                                                                     //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_startofpacket  (1'b0),                                                                            // (terminated)
		.in_endofpacket    (1'b0),                                                                            // (terminated)
		.out_startofpacket (),                                                                                // (terminated)
		.out_endofpacket   (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_BEGIN_BURST           (63),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.PKT_BURST_TYPE_H          (60),
		.PKT_BURST_TYPE_L          (59),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_TRANS_EXCLUSIVE       (51),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_THREAD_ID_H           (73),
		.PKT_THREAD_ID_L           (73),
		.PKT_CACHE_H               (80),
		.PKT_CACHE_L               (77),
		.PKT_DATA_SIDEBAND_H       (62),
		.PKT_DATA_SIDEBAND_L       (62),
		.PKT_QOS_H                 (64),
		.PKT_QOS_L                 (64),
		.PKT_ADDR_SIDEBAND_H       (61),
		.PKT_ADDR_SIDEBAND_L       (61),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.ST_DATA_W                 (83),
		.ST_CHANNEL_W              (11),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (1),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) apb_m0_translator_avalon_universal_master_0_agent (
		.clk                     (syspll_c0_clk),                                                      //       clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                 // clk_reset.reset
		.av_address              (apb_m0_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (apb_m0_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (apb_m0_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (apb_m0_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (apb_m0_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (apb_m0_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (apb_m0_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (apb_m0_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (apb_m0_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (apb_m0_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (apb_m0_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (apb_m0_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (apb_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (apb_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (apb_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (apb_m0_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (limiter_001_rsp_src_valid),                                          //        rp.valid
		.rp_data                 (limiter_001_rsp_src_data),                                           //          .data
		.rp_channel              (limiter_001_rsp_src_channel),                                        //          .channel
		.rp_startofpacket        (limiter_001_rsp_src_startofpacket),                                  //          .startofpacket
		.rp_endofpacket          (limiter_001_rsp_src_endofpacket),                                    //          .endofpacket
		.rp_ready                (limiter_001_rsp_src_ready),                                          //          .ready
		.av_response             (),                                                                   // (terminated)
		.av_writeresponserequest (1'b0),                                                               // (terminated)
		.av_writeresponsevalid   ()                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (syspll_c0_clk),                                                                                    //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                               //       clk_reset.reset
		.m0_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_004_src0_ready),                                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_004_src0_valid),                                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_004_src0_data),                                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_004_src0_startofpacket),                                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_004_src0_endofpacket),                                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_004_src0_channel),                                                                  //                .channel
		.rf_sink_ready           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (syspll_c0_clk),                                                                                    //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                               // clk_reset.reset
		.in_data           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                             // (terminated)
		.almost_full_data  (),                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                             // (terminated)
		.out_empty         (),                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                             // (terminated)
		.out_error         (),                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                             // (terminated)
		.out_channel       ()                                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) timer_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (syspll_c0_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                            //       clk_reset.reset
		.m0_address              (timer_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_004_src1_ready),                                                 //              cp.ready
		.cp_valid                (cmd_xbar_demux_004_src1_valid),                                                 //                .valid
		.cp_data                 (cmd_xbar_demux_004_src1_data),                                                  //                .data
		.cp_startofpacket        (cmd_xbar_demux_004_src1_startofpacket),                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_004_src1_endofpacket),                                           //                .endofpacket
		.cp_channel              (cmd_xbar_demux_004_src1_channel),                                               //                .channel
		.rf_sink_ready           (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (syspll_c0_clk),                                                                 //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                            // clk_reset.reset
		.in_data           (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) uart0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (syspll_c0_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                            //       clk_reset.reset
		.m0_address              (uart0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (uart0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (uart0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (uart0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (uart0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (uart0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (uart0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (uart0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (uart0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (uart0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (uart0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (uart0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (uart0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (uart0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (uart0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (uart0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_004_src2_ready),                                                 //              cp.ready
		.cp_valid                (cmd_xbar_demux_004_src2_valid),                                                 //                .valid
		.cp_data                 (cmd_xbar_demux_004_src2_data),                                                  //                .data
		.cp_startofpacket        (cmd_xbar_demux_004_src2_startofpacket),                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_004_src2_endofpacket),                                           //                .endofpacket
		.cp_channel              (cmd_xbar_demux_004_src2_channel),                                               //                .channel
		.rf_sink_ready           (uart0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (uart0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (uart0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (uart0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (uart0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (uart0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (uart0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (uart0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (uart0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (uart0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (uart0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (uart0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (uart0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (uart0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (uart0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (uart0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) uart0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (syspll_c0_clk),                                                                 //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                            // clk_reset.reset
		.in_data           (uart0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (uart0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (uart0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (uart0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (uart0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (uart0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (uart0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (uart0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (uart0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (uart0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sw_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (syspll_c0_clk),                                                              //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                         //       clk_reset.reset
		.m0_address              (sw_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sw_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sw_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sw_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sw_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sw_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sw_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sw_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sw_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sw_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sw_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sw_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sw_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sw_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sw_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sw_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_004_src3_ready),                                              //              cp.ready
		.cp_valid                (cmd_xbar_demux_004_src3_valid),                                              //                .valid
		.cp_data                 (cmd_xbar_demux_004_src3_data),                                               //                .data
		.cp_startofpacket        (cmd_xbar_demux_004_src3_startofpacket),                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_004_src3_endofpacket),                                        //                .endofpacket
		.cp_channel              (cmd_xbar_demux_004_src3_channel),                                            //                .channel
		.rf_sink_ready           (sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sw_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sw_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sw_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sw_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sw_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                      //     (terminated)
		.m0_writeresponserequest (),                                                                           //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                        //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (syspll_c0_clk),                                                              //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                         // clk_reset.reset
		.in_data           (sw_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sw_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sw_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sw_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sw_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                      // (terminated)
		.csr_read          (1'b0),                                                                       // (terminated)
		.csr_write         (1'b0),                                                                       // (terminated)
		.csr_readdata      (),                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                       // (terminated)
		.almost_full_data  (),                                                                           // (terminated)
		.almost_empty_data (),                                                                           // (terminated)
		.in_empty          (1'b0),                                                                       // (terminated)
		.out_empty         (),                                                                           // (terminated)
		.in_error          (1'b0),                                                                       // (terminated)
		.out_error         (),                                                                           // (terminated)
		.in_channel        (1'b0),                                                                       // (terminated)
		.out_channel       ()                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) led_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (syspll_c0_clk),                                                               //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                          //       clk_reset.reset
		.m0_address              (led_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (led_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (led_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (led_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (led_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (led_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (led_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (led_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (led_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (led_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (led_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (led_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (led_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (led_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (led_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (led_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_004_src4_ready),                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_004_src4_valid),                                               //                .valid
		.cp_data                 (cmd_xbar_demux_004_src4_data),                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_004_src4_startofpacket),                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_004_src4_endofpacket),                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_004_src4_channel),                                             //                .channel
		.rf_sink_ready           (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (led_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (led_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (led_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (led_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (led_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                       //     (terminated)
		.m0_writeresponserequest (),                                                                            //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                         //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (syspll_c0_clk),                                                               //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.in_data           (led_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (led_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (led_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (led_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (led_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                       // (terminated)
		.csr_read          (1'b0),                                                                        // (terminated)
		.csr_write         (1'b0),                                                                        // (terminated)
		.csr_readdata      (),                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                        // (terminated)
		.almost_full_data  (),                                                                            // (terminated)
		.almost_empty_data (),                                                                            // (terminated)
		.in_empty          (1'b0),                                                                        // (terminated)
		.out_empty         (),                                                                            // (terminated)
		.in_error          (1'b0),                                                                        // (terminated)
		.out_error         (),                                                                            // (terminated)
		.in_channel        (1'b0),                                                                        // (terminated)
		.out_channel       ()                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) button1_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (syspll_c0_clk),                                                                   //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (button1_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (button1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (button1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (button1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (button1_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (button1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (button1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (button1_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (button1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (button1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (button1_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (button1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (button1_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (button1_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (button1_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (button1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_004_src5_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_004_src5_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_004_src5_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_004_src5_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_004_src5_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_004_src5_channel),                                                 //                .channel
		.rf_sink_ready           (button1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (button1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (button1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (button1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (button1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (button1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (button1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (button1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (button1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (button1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (button1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (button1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (button1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (button1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (button1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (button1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) button1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (syspll_c0_clk),                                                                   //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                              // clk_reset.reset
		.in_data           (button1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (button1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (button1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (button1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (button1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (button1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (button1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (button1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (button1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (button1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) button2_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (syspll_c0_clk),                                                                   //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (button2_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (button2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (button2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (button2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (button2_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (button2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (button2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (button2_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (button2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (button2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (button2_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (button2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (button2_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (button2_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (button2_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (button2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_004_src6_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_004_src6_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_004_src6_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_004_src6_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_004_src6_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_004_src6_channel),                                                 //                .channel
		.rf_sink_ready           (button2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (button2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (button2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (button2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (button2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (button2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (button2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (button2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (button2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (button2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (button2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (button2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (button2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (button2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (button2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (button2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) button2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (syspll_c0_clk),                                                                   //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                              // clk_reset.reset
		.in_data           (button2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (button2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (button2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (button2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (button2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (button2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (button2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (button2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (button2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (button2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) hex0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (syspll_c0_clk),                                                                //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                           //       clk_reset.reset
		.m0_address              (hex0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (hex0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (hex0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (hex0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (hex0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (hex0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (hex0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (hex0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (hex0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (hex0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (hex0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (hex0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (hex0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (hex0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (hex0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (hex0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_004_src7_ready),                                                //              cp.ready
		.cp_valid                (cmd_xbar_demux_004_src7_valid),                                                //                .valid
		.cp_data                 (cmd_xbar_demux_004_src7_data),                                                 //                .data
		.cp_startofpacket        (cmd_xbar_demux_004_src7_startofpacket),                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_004_src7_endofpacket),                                          //                .endofpacket
		.cp_channel              (cmd_xbar_demux_004_src7_channel),                                              //                .channel
		.rf_sink_ready           (hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (hex0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (hex0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (hex0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (hex0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (hex0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (hex0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (syspll_c0_clk),                                                                //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.in_data           (hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) hex1_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (syspll_c0_clk),                                                                //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                           //       clk_reset.reset
		.m0_address              (hex1_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (hex1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (hex1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (hex1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (hex1_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (hex1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (hex1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (hex1_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (hex1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (hex1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (hex1_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (hex1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (hex1_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (hex1_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (hex1_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (hex1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_004_src8_ready),                                                //              cp.ready
		.cp_valid                (cmd_xbar_demux_004_src8_valid),                                                //                .valid
		.cp_data                 (cmd_xbar_demux_004_src8_data),                                                 //                .data
		.cp_startofpacket        (cmd_xbar_demux_004_src8_startofpacket),                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_004_src8_endofpacket),                                          //                .endofpacket
		.cp_channel              (cmd_xbar_demux_004_src8_channel),                                              //                .channel
		.rf_sink_ready           (hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (hex1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (hex1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (hex1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (hex1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (hex1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (hex1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (syspll_c0_clk),                                                                //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.in_data           (hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) hex2_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (syspll_c0_clk),                                                                //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                           //       clk_reset.reset
		.m0_address              (hex2_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (hex2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (hex2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (hex2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (hex2_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (hex2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (hex2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (hex2_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (hex2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (hex2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (hex2_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (hex2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (hex2_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (hex2_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (hex2_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (hex2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_004_src9_ready),                                                //              cp.ready
		.cp_valid                (cmd_xbar_demux_004_src9_valid),                                                //                .valid
		.cp_data                 (cmd_xbar_demux_004_src9_data),                                                 //                .data
		.cp_startofpacket        (cmd_xbar_demux_004_src9_startofpacket),                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_004_src9_endofpacket),                                          //                .endofpacket
		.cp_channel              (cmd_xbar_demux_004_src9_channel),                                              //                .channel
		.rf_sink_ready           (hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (hex2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (hex2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (hex2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (hex2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (hex2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (hex2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (syspll_c0_clk),                                                                //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.in_data           (hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) hex3_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (syspll_c0_clk),                                                                //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                           //       clk_reset.reset
		.m0_address              (hex3_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (hex3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (hex3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (hex3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (hex3_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (hex3_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (hex3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (hex3_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (hex3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (hex3_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (hex3_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (hex3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (hex3_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (hex3_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (hex3_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (hex3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_004_src10_ready),                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_004_src10_valid),                                               //                .valid
		.cp_data                 (cmd_xbar_demux_004_src10_data),                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_004_src10_startofpacket),                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_004_src10_endofpacket),                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_004_src10_channel),                                             //                .channel
		.rf_sink_ready           (hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (hex3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (hex3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (hex3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (hex3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (hex3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (hex3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (syspll_c0_clk),                                                                //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.in_data           (hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	DE0Qsys_addr_router addr_router (
		.sink_ready         (nios2cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (syspll_c0_clk),                                                                           //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                      // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                   //       src.ready
		.src_valid          (addr_router_src_valid),                                                                   //          .valid
		.src_data           (addr_router_src_data),                                                                    //          .data
		.src_channel        (addr_router_src_channel),                                                                 //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                           //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                              //          .endofpacket
	);

	DE0Qsys_addr_router_001 addr_router_001 (
		.sink_ready         (dma_write_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (dma_write_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (dma_write_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (dma_write_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (dma_write_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (syspll_c0_clk),                                                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                    //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                    //          .valid
		.src_data           (addr_router_001_src_data),                                                     //          .data
		.src_channel        (addr_router_001_src_channel),                                                  //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                               //          .endofpacket
	);

	DE0Qsys_addr_router_002 addr_router_002 (
		.sink_ready         (nios2cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2cpu_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (syspll_c0_clk),                                                                    //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (addr_router_002_src_ready),                                                        //       src.ready
		.src_valid          (addr_router_002_src_valid),                                                        //          .valid
		.src_data           (addr_router_002_src_data),                                                         //          .data
		.src_channel        (addr_router_002_src_channel),                                                      //          .channel
		.src_startofpacket  (addr_router_002_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (addr_router_002_src_endofpacket)                                                   //          .endofpacket
	);

	DE0Qsys_addr_router_001 addr_router_003 (
		.sink_ready         (dma_read_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (dma_read_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (dma_read_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (dma_read_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (dma_read_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (syspll_c0_clk),                                                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (addr_router_003_src_ready),                                                   //       src.ready
		.src_valid          (addr_router_003_src_valid),                                                   //          .valid
		.src_data           (addr_router_003_src_data),                                                    //          .data
		.src_channel        (addr_router_003_src_channel),                                                 //          .channel
		.src_startofpacket  (addr_router_003_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (addr_router_003_src_endofpacket)                                              //          .endofpacket
	);

	DE0Qsys_id_router id_router (
		.sink_ready         (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (syspll_c0_clk),                                                                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                   //       src.ready
		.src_valid          (id_router_src_valid),                                                                   //          .valid
		.src_data           (id_router_src_data),                                                                    //          .data
		.src_channel        (id_router_src_channel),                                                                 //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                           //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                              //          .endofpacket
	);

	DE0Qsys_id_router_001 id_router_001 (
		.sink_ready         (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (syspll_c0_clk),                                                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                  //       src.ready
		.src_valid          (id_router_001_src_valid),                                                  //          .valid
		.src_data           (id_router_001_src_data),                                                   //          .data
		.src_channel        (id_router_001_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                             //          .endofpacket
	);

	DE0Qsys_id_router id_router_002 (
		.sink_ready         (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (syspll_c0_clk),                                                                     //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                           //       src.ready
		.src_valid          (id_router_002_src_valid),                                                           //          .valid
		.src_data           (id_router_002_src_data),                                                            //          .data
		.src_channel        (id_router_002_src_channel),                                                         //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                                   //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                                      //          .endofpacket
	);

	DE0Qsys_id_router_003 id_router_003 (
		.sink_ready         (apb_s0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (apb_s0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (apb_s0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (apb_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (apb_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (syspll_c0_clk),                                                     //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                           //       src.ready
		.src_valid          (id_router_003_src_valid),                                           //          .valid
		.src_data           (id_router_003_src_data),                                            //          .data
		.src_channel        (id_router_003_src_channel),                                         //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                   //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                      //          .endofpacket
	);

	DE0Qsys_id_router_004 id_router_004 (
		.sink_ready         (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_50m_clk),                                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                     //       src.ready
		.src_valid          (id_router_004_src_valid),                                                     //          .valid
		.src_data           (id_router_004_src_data),                                                      //          .data
		.src_channel        (id_router_004_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                                //          .endofpacket
	);

	DE0Qsys_addr_router_004 addr_router_004 (
		.sink_ready         (apb_m0_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (apb_m0_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (apb_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (apb_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (apb_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (syspll_c0_clk),                                                      //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                 // clk_reset.reset
		.src_ready          (addr_router_004_src_ready),                                          //       src.ready
		.src_valid          (addr_router_004_src_valid),                                          //          .valid
		.src_data           (addr_router_004_src_data),                                           //          .data
		.src_channel        (addr_router_004_src_channel),                                        //          .channel
		.src_startofpacket  (addr_router_004_src_startofpacket),                                  //          .startofpacket
		.src_endofpacket    (addr_router_004_src_endofpacket)                                     //          .endofpacket
	);

	DE0Qsys_id_router_005 id_router_005 (
		.sink_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (syspll_c0_clk),                                                                          //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                                //       src.ready
		.src_valid          (id_router_005_src_valid),                                                                //          .valid
		.src_data           (id_router_005_src_data),                                                                 //          .data
		.src_channel        (id_router_005_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                                           //          .endofpacket
	);

	DE0Qsys_id_router_005 id_router_006 (
		.sink_ready         (timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (syspll_c0_clk),                                                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                  // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                             //       src.ready
		.src_valid          (id_router_006_src_valid),                                             //          .valid
		.src_data           (id_router_006_src_data),                                              //          .data
		.src_channel        (id_router_006_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                        //          .endofpacket
	);

	DE0Qsys_id_router_005 id_router_007 (
		.sink_ready         (uart0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (uart0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (uart0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (uart0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (uart0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (syspll_c0_clk),                                                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                  // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                             //       src.ready
		.src_valid          (id_router_007_src_valid),                                             //          .valid
		.src_data           (id_router_007_src_data),                                              //          .data
		.src_channel        (id_router_007_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                        //          .endofpacket
	);

	DE0Qsys_id_router_005 id_router_008 (
		.sink_ready         (sw_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sw_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sw_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sw_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sw_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (syspll_c0_clk),                                                    //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                               // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                          //       src.ready
		.src_valid          (id_router_008_src_valid),                                          //          .valid
		.src_data           (id_router_008_src_data),                                           //          .data
		.src_channel        (id_router_008_src_channel),                                        //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                  //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                     //          .endofpacket
	);

	DE0Qsys_id_router_005 id_router_009 (
		.sink_ready         (led_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (led_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (led_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (led_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (led_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (syspll_c0_clk),                                                     //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                           //       src.ready
		.src_valid          (id_router_009_src_valid),                                           //          .valid
		.src_data           (id_router_009_src_data),                                            //          .data
		.src_channel        (id_router_009_src_channel),                                         //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                   //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                      //          .endofpacket
	);

	DE0Qsys_id_router_005 id_router_010 (
		.sink_ready         (button1_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (button1_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (button1_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (button1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (button1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (syspll_c0_clk),                                                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                               //       src.ready
		.src_valid          (id_router_010_src_valid),                                               //          .valid
		.src_data           (id_router_010_src_data),                                                //          .data
		.src_channel        (id_router_010_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                          //          .endofpacket
	);

	DE0Qsys_id_router_005 id_router_011 (
		.sink_ready         (button2_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (button2_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (button2_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (button2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (button2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (syspll_c0_clk),                                                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_011_src_ready),                                               //       src.ready
		.src_valid          (id_router_011_src_valid),                                               //          .valid
		.src_data           (id_router_011_src_data),                                                //          .data
		.src_channel        (id_router_011_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_011_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_011_src_endofpacket)                                          //          .endofpacket
	);

	DE0Qsys_id_router_005 id_router_012 (
		.sink_ready         (hex0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (hex0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (hex0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (hex0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (hex0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (syspll_c0_clk),                                                      //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                 // clk_reset.reset
		.src_ready          (id_router_012_src_ready),                                            //       src.ready
		.src_valid          (id_router_012_src_valid),                                            //          .valid
		.src_data           (id_router_012_src_data),                                             //          .data
		.src_channel        (id_router_012_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_012_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_012_src_endofpacket)                                       //          .endofpacket
	);

	DE0Qsys_id_router_005 id_router_013 (
		.sink_ready         (hex1_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (hex1_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (hex1_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (hex1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (hex1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (syspll_c0_clk),                                                      //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                 // clk_reset.reset
		.src_ready          (id_router_013_src_ready),                                            //       src.ready
		.src_valid          (id_router_013_src_valid),                                            //          .valid
		.src_data           (id_router_013_src_data),                                             //          .data
		.src_channel        (id_router_013_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_013_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_013_src_endofpacket)                                       //          .endofpacket
	);

	DE0Qsys_id_router_005 id_router_014 (
		.sink_ready         (hex2_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (hex2_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (hex2_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (hex2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (hex2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (syspll_c0_clk),                                                      //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                 // clk_reset.reset
		.src_ready          (id_router_014_src_ready),                                            //       src.ready
		.src_valid          (id_router_014_src_valid),                                            //          .valid
		.src_data           (id_router_014_src_data),                                             //          .data
		.src_channel        (id_router_014_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_014_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_014_src_endofpacket)                                       //          .endofpacket
	);

	DE0Qsys_id_router_005 id_router_015 (
		.sink_ready         (hex3_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (hex3_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (hex3_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (hex3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (hex3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (syspll_c0_clk),                                                      //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                 // clk_reset.reset
		.src_ready          (id_router_015_src_ready),                                            //       src.ready
		.src_valid          (id_router_015_src_valid),                                            //          .valid
		.src_data           (id_router_015_src_data),                                             //          .data
		.src_channel        (id_router_015_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_015_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_015_src_endofpacket)                                       //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (95),
		.PKT_DEST_ID_L             (93),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.MAX_OUTSTANDING_RESPONSES (9),
		.PIPELINED                 (0),
		.ST_DATA_W                 (106),
		.ST_CHANNEL_W              (5),
		.VALID_WIDTH               (5),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (77),
		.PKT_BYTE_CNT_L            (68),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (syspll_c0_clk),                      //       clk.clk
		.reset                  (rst_controller_001_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_003_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_003_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_003_src_data),           //          .data
		.cmd_sink_channel       (addr_router_003_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_003_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_003_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),              //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),               //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),            //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),      //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),        //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_003_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_003_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_003_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_003_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_003_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_003_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),              //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),              //          .valid
		.rsp_src_data           (limiter_rsp_src_data),               //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),            //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),      //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),        //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)              // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.MAX_OUTSTANDING_RESPONSES (1),
		.PIPELINED                 (0),
		.ST_DATA_W                 (83),
		.ST_CHANNEL_W              (11),
		.VALID_WIDTH               (11),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_001 (
		.clk                    (syspll_c0_clk),                      //       clk.clk
		.reset                  (rst_controller_001_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_004_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_004_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_004_src_data),           //          .data
		.cmd_sink_channel       (addr_router_004_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_004_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_004_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_001_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_001_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_001_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_001_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_001_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_004_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_004_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_004_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_004_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_004_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_004_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_001_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_001_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_001_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_001_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_001_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_001_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_001_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (43),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (70),
		.PKT_BYTE_CNT_H            (59),
		.PKT_BYTE_CNT_L            (50),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURST_SIZE_H          (65),
		.PKT_BURST_SIZE_L          (63),
		.PKT_BURST_TYPE_H          (67),
		.PKT_BURST_TYPE_L          (66),
		.PKT_BURSTWRAP_H           (62),
		.PKT_BURSTWRAP_L           (60),
		.PKT_TRANS_COMPRESSED_READ (44),
		.PKT_TRANS_WRITE           (46),
		.PKT_TRANS_READ            (47),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (88),
		.ST_CHANNEL_W              (5),
		.OUT_BYTE_CNT_H            (51),
		.OUT_BURSTWRAP_H           (62),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter (
		.clk                   (syspll_c0_clk),                       //       cr0.clk
		.reset                 (rst_controller_001_reset_out_reset),  // cr0_reset.reset
		.sink0_valid           (width_adapter_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_src_data),              //          .data
		.sink0_channel         (width_adapter_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_src_ready),             //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (88),
		.PKT_BYTE_CNT_H            (77),
		.PKT_BYTE_CNT_L            (68),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (83),
		.PKT_BURST_SIZE_L          (81),
		.PKT_BURST_TYPE_H          (85),
		.PKT_BURST_TYPE_L          (84),
		.PKT_BURSTWRAP_H           (80),
		.PKT_BURSTWRAP_L           (78),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (106),
		.ST_CHANNEL_W              (5),
		.OUT_BYTE_CNT_H            (70),
		.OUT_BURSTWRAP_H           (80),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter_001 (
		.clk                   (syspll_c0_clk),                           //       cr0.clk
		.reset                 (rst_controller_001_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (cmd_xbar_mux_003_src_valid),              //     sink0.valid
		.sink0_data            (cmd_xbar_mux_003_src_data),               //          .data
		.sink0_channel         (cmd_xbar_mux_003_src_channel),            //          .channel
		.sink0_startofpacket   (cmd_xbar_mux_003_src_startofpacket),      //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_mux_003_src_endofpacket),        //          .endofpacket
		.sink0_ready           (cmd_xbar_mux_003_src_ready),              //          .ready
		.source0_valid         (burst_adapter_001_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_001_source0_data),          //          .data
		.source0_channel       (burst_adapter_001_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_001_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_001_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_001_source0_ready)          //          .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                 // reset_in0.reset
		.clk        (clk_50m_clk),                    //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req  (),                               // (terminated)
		.reset_in1  (1'b0),                           // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_001 (
		.reset_in0  (~reset_reset_n),                         // reset_in0.reset
		.reset_in1  (nios2cpu_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (syspll_c0_clk),                          //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req  (),                                       // (terminated)
		.reset_in2  (1'b0),                                   // (terminated)
		.reset_in3  (1'b0),                                   // (terminated)
		.reset_in4  (1'b0),                                   // (terminated)
		.reset_in5  (1'b0),                                   // (terminated)
		.reset_in6  (1'b0),                                   // (terminated)
		.reset_in7  (1'b0),                                   // (terminated)
		.reset_in8  (1'b0),                                   // (terminated)
		.reset_in9  (1'b0),                                   // (terminated)
		.reset_in10 (1'b0),                                   // (terminated)
		.reset_in11 (1'b0),                                   // (terminated)
		.reset_in12 (1'b0),                                   // (terminated)
		.reset_in13 (1'b0),                                   // (terminated)
		.reset_in14 (1'b0),                                   // (terminated)
		.reset_in15 (1'b0)                                    // (terminated)
	);

	DE0Qsys_cmd_xbar_demux cmd_xbar_demux (
		.clk                (syspll_c0_clk),                      //       clk.clk
		.reset              (rst_controller_001_reset_out_reset), // clk_reset.reset
		.sink_ready         (addr_router_src_ready),              //      sink.ready
		.sink_channel       (addr_router_src_channel),            //          .channel
		.sink_data          (addr_router_src_data),               //          .data
		.sink_startofpacket (addr_router_src_startofpacket),      //          .startofpacket
		.sink_endofpacket   (addr_router_src_endofpacket),        //          .endofpacket
		.sink_valid         (addr_router_src_valid),              //          .valid
		.src0_ready         (cmd_xbar_demux_src0_ready),          //      src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),          //          .valid
		.src0_data          (cmd_xbar_demux_src0_data),           //          .data
		.src0_channel       (cmd_xbar_demux_src0_channel),        //          .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),    //          .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),          //      src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),          //          .valid
		.src1_data          (cmd_xbar_demux_src1_data),           //          .data
		.src1_channel       (cmd_xbar_demux_src1_channel),        //          .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),    //          .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),          //      src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),          //          .valid
		.src2_data          (cmd_xbar_demux_src2_data),           //          .data
		.src2_channel       (cmd_xbar_demux_src2_channel),        //          .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket),  //          .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket),    //          .endofpacket
		.src3_ready         (cmd_xbar_demux_src3_ready),          //      src3.ready
		.src3_valid         (cmd_xbar_demux_src3_valid),          //          .valid
		.src3_data          (cmd_xbar_demux_src3_data),           //          .data
		.src3_channel       (cmd_xbar_demux_src3_channel),        //          .channel
		.src3_startofpacket (cmd_xbar_demux_src3_startofpacket),  //          .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_src3_endofpacket)     //          .endofpacket
	);

	DE0Qsys_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                (syspll_c0_clk),                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_001_src_ready),             //      sink.ready
		.sink_channel       (addr_router_001_src_channel),           //          .channel
		.sink_data          (addr_router_001_src_data),              //          .data
		.sink_startofpacket (addr_router_001_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_001_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_001_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	DE0Qsys_cmd_xbar_demux_002 cmd_xbar_demux_002 (
		.clk                (syspll_c0_clk),                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_002_src_ready),             //      sink.ready
		.sink_channel       (addr_router_002_src_channel),           //          .channel
		.sink_data          (addr_router_002_src_data),              //          .data
		.sink_startofpacket (addr_router_002_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_002_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_002_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.src2_ready         (cmd_xbar_demux_002_src2_ready),         //      src2.ready
		.src2_valid         (cmd_xbar_demux_002_src2_valid),         //          .valid
		.src2_data          (cmd_xbar_demux_002_src2_data),          //          .data
		.src2_channel       (cmd_xbar_demux_002_src2_channel),       //          .channel
		.src2_startofpacket (cmd_xbar_demux_002_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_002_src2_endofpacket),   //          .endofpacket
		.src3_ready         (cmd_xbar_demux_002_src3_ready),         //      src3.ready
		.src3_valid         (cmd_xbar_demux_002_src3_valid),         //          .valid
		.src3_data          (cmd_xbar_demux_002_src3_data),          //          .data
		.src3_channel       (cmd_xbar_demux_002_src3_channel),       //          .channel
		.src3_startofpacket (cmd_xbar_demux_002_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_002_src3_endofpacket),   //          .endofpacket
		.src4_ready         (cmd_xbar_demux_002_src4_ready),         //      src4.ready
		.src4_valid         (cmd_xbar_demux_002_src4_valid),         //          .valid
		.src4_data          (cmd_xbar_demux_002_src4_data),          //          .data
		.src4_channel       (cmd_xbar_demux_002_src4_channel),       //          .channel
		.src4_startofpacket (cmd_xbar_demux_002_src4_startofpacket), //          .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_002_src4_endofpacket)    //          .endofpacket
	);

	DE0Qsys_cmd_xbar_demux_003 cmd_xbar_demux_003 (
		.clk                (syspll_c0_clk),                         //        clk.clk
		.reset              (rst_controller_001_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),                 //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),               //           .channel
		.sink_data          (limiter_cmd_src_data),                  //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),         //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),           //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),                // sink_valid.data
		.src0_ready         (cmd_xbar_demux_003_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_003_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_003_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_003_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_003_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_003_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_003_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_003_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_003_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_003_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_003_src1_endofpacket)    //           .endofpacket
	);

	DE0Qsys_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (syspll_c0_clk),                         //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	DE0Qsys_cmd_xbar_mux_001 cmd_xbar_mux_001 (
		.clk                 (syspll_c0_clk),                         //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_002_src1_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_002_src1_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_002_src1_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_002_src1_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	DE0Qsys_cmd_xbar_mux cmd_xbar_mux_002 (
		.clk                 (syspll_c0_clk),                         //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_002_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_002_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src2_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src2_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src2_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src2_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src2_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src2_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_002_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src2_endofpacket)    //          .endofpacket
	);

	DE0Qsys_cmd_xbar_mux_001 cmd_xbar_mux_003 (
		.clk                 (syspll_c0_clk),                         //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_003_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_003_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_003_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_003_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_003_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_003_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src3_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src3_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src3_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src3_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src3_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src3_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_002_src3_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_002_src3_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_002_src3_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_002_src3_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_002_src3_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_002_src3_endofpacket),   //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_003_src1_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_003_src1_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_003_src1_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_003_src1_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_003_src1_endofpacket)    //          .endofpacket
	);

	DE0Qsys_cmd_xbar_demux_001 rsp_xbar_demux (
		.clk                (syspll_c0_clk),                      //       clk.clk
		.reset              (rst_controller_001_reset_out_reset), // clk_reset.reset
		.sink_ready         (id_router_src_ready),                //      sink.ready
		.sink_channel       (id_router_src_channel),              //          .channel
		.sink_data          (id_router_src_data),                 //          .data
		.sink_startofpacket (id_router_src_startofpacket),        //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),          //          .endofpacket
		.sink_valid         (id_router_src_valid),                //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),          //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),          //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),           //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),        //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),    //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),          //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),          //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),           //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),        //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)     //          .endofpacket
	);

	DE0Qsys_cmd_xbar_demux rsp_xbar_demux_001 (
		.clk                (syspll_c0_clk),                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (width_adapter_001_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_001_src_channel),         //          .channel
		.sink_data          (width_adapter_001_src_data),            //          .data
		.sink_startofpacket (width_adapter_001_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_001_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_001_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_001_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_001_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_001_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_001_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_001_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_001_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_001_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_001_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_001_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_001_src3_endofpacket)    //          .endofpacket
	);

	DE0Qsys_cmd_xbar_demux_001 rsp_xbar_demux_002 (
		.clk                (syspll_c0_clk),                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket)    //          .endofpacket
	);

	DE0Qsys_cmd_xbar_demux rsp_xbar_demux_003 (
		.clk                (syspll_c0_clk),                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_003_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_003_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_003_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_003_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_003_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_003_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_003_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_003_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_003_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_003_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_003_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_003_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_003_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_003_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_003_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_003_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_003_src3_endofpacket)    //          .endofpacket
	);

	DE0Qsys_rsp_xbar_demux_004 rsp_xbar_demux_004 (
		.clk                (clk_50m_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	DE0Qsys_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (syspll_c0_clk),                         //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	DE0Qsys_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                 (syspll_c0_clk),                         //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_001_src1_ready),         //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink0_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink0_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.sink0_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_003_src1_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_003_src1_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_003_src1_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_003_src1_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_003_src1_endofpacket)    //          .endofpacket
	);

	DE0Qsys_rsp_xbar_mux_002 rsp_xbar_mux_002 (
		.clk                 (syspll_c0_clk),                         //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_002_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_002_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src2_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src2_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src2_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src2_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src2_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src1_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src2_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src2_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src2_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_003_src2_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src2_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src2_endofpacket),   //          .endofpacket
		.sink4_ready         (crosser_001_out_ready),                 //     sink4.ready
		.sink4_valid         (crosser_001_out_valid),                 //          .valid
		.sink4_channel       (crosser_001_out_channel),               //          .channel
		.sink4_data          (crosser_001_out_data),                  //          .data
		.sink4_startofpacket (crosser_001_out_startofpacket),         //          .startofpacket
		.sink4_endofpacket   (crosser_001_out_endofpacket)            //          .endofpacket
	);

	DE0Qsys_rsp_xbar_mux_001 rsp_xbar_mux_003 (
		.clk                 (syspll_c0_clk),                         //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_003_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_003_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_003_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_003_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_003_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_003_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_001_src3_ready),         //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_001_src3_valid),         //          .valid
		.sink0_channel       (rsp_xbar_demux_001_src3_channel),       //          .channel
		.sink0_data          (rsp_xbar_demux_001_src3_data),          //          .data
		.sink0_startofpacket (rsp_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_001_src3_endofpacket),   //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_003_src3_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_003_src3_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_003_src3_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_003_src3_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_003_src3_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_003_src3_endofpacket)    //          .endofpacket
	);

	DE0Qsys_cmd_xbar_demux_004 cmd_xbar_demux_004 (
		.clk                 (syspll_c0_clk),                          //        clk.clk
		.reset               (rst_controller_001_reset_out_reset),     //  clk_reset.reset
		.sink_ready          (limiter_001_cmd_src_ready),              //       sink.ready
		.sink_channel        (limiter_001_cmd_src_channel),            //           .channel
		.sink_data           (limiter_001_cmd_src_data),               //           .data
		.sink_startofpacket  (limiter_001_cmd_src_startofpacket),      //           .startofpacket
		.sink_endofpacket    (limiter_001_cmd_src_endofpacket),        //           .endofpacket
		.sink_valid          (limiter_001_cmd_valid_data),             // sink_valid.data
		.src0_ready          (cmd_xbar_demux_004_src0_ready),          //       src0.ready
		.src0_valid          (cmd_xbar_demux_004_src0_valid),          //           .valid
		.src0_data           (cmd_xbar_demux_004_src0_data),           //           .data
		.src0_channel        (cmd_xbar_demux_004_src0_channel),        //           .channel
		.src0_startofpacket  (cmd_xbar_demux_004_src0_startofpacket),  //           .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_004_src0_endofpacket),    //           .endofpacket
		.src1_ready          (cmd_xbar_demux_004_src1_ready),          //       src1.ready
		.src1_valid          (cmd_xbar_demux_004_src1_valid),          //           .valid
		.src1_data           (cmd_xbar_demux_004_src1_data),           //           .data
		.src1_channel        (cmd_xbar_demux_004_src1_channel),        //           .channel
		.src1_startofpacket  (cmd_xbar_demux_004_src1_startofpacket),  //           .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_004_src1_endofpacket),    //           .endofpacket
		.src2_ready          (cmd_xbar_demux_004_src2_ready),          //       src2.ready
		.src2_valid          (cmd_xbar_demux_004_src2_valid),          //           .valid
		.src2_data           (cmd_xbar_demux_004_src2_data),           //           .data
		.src2_channel        (cmd_xbar_demux_004_src2_channel),        //           .channel
		.src2_startofpacket  (cmd_xbar_demux_004_src2_startofpacket),  //           .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_004_src2_endofpacket),    //           .endofpacket
		.src3_ready          (cmd_xbar_demux_004_src3_ready),          //       src3.ready
		.src3_valid          (cmd_xbar_demux_004_src3_valid),          //           .valid
		.src3_data           (cmd_xbar_demux_004_src3_data),           //           .data
		.src3_channel        (cmd_xbar_demux_004_src3_channel),        //           .channel
		.src3_startofpacket  (cmd_xbar_demux_004_src3_startofpacket),  //           .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_004_src3_endofpacket),    //           .endofpacket
		.src4_ready          (cmd_xbar_demux_004_src4_ready),          //       src4.ready
		.src4_valid          (cmd_xbar_demux_004_src4_valid),          //           .valid
		.src4_data           (cmd_xbar_demux_004_src4_data),           //           .data
		.src4_channel        (cmd_xbar_demux_004_src4_channel),        //           .channel
		.src4_startofpacket  (cmd_xbar_demux_004_src4_startofpacket),  //           .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_004_src4_endofpacket),    //           .endofpacket
		.src5_ready          (cmd_xbar_demux_004_src5_ready),          //       src5.ready
		.src5_valid          (cmd_xbar_demux_004_src5_valid),          //           .valid
		.src5_data           (cmd_xbar_demux_004_src5_data),           //           .data
		.src5_channel        (cmd_xbar_demux_004_src5_channel),        //           .channel
		.src5_startofpacket  (cmd_xbar_demux_004_src5_startofpacket),  //           .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_004_src5_endofpacket),    //           .endofpacket
		.src6_ready          (cmd_xbar_demux_004_src6_ready),          //       src6.ready
		.src6_valid          (cmd_xbar_demux_004_src6_valid),          //           .valid
		.src6_data           (cmd_xbar_demux_004_src6_data),           //           .data
		.src6_channel        (cmd_xbar_demux_004_src6_channel),        //           .channel
		.src6_startofpacket  (cmd_xbar_demux_004_src6_startofpacket),  //           .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_004_src6_endofpacket),    //           .endofpacket
		.src7_ready          (cmd_xbar_demux_004_src7_ready),          //       src7.ready
		.src7_valid          (cmd_xbar_demux_004_src7_valid),          //           .valid
		.src7_data           (cmd_xbar_demux_004_src7_data),           //           .data
		.src7_channel        (cmd_xbar_demux_004_src7_channel),        //           .channel
		.src7_startofpacket  (cmd_xbar_demux_004_src7_startofpacket),  //           .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_004_src7_endofpacket),    //           .endofpacket
		.src8_ready          (cmd_xbar_demux_004_src8_ready),          //       src8.ready
		.src8_valid          (cmd_xbar_demux_004_src8_valid),          //           .valid
		.src8_data           (cmd_xbar_demux_004_src8_data),           //           .data
		.src8_channel        (cmd_xbar_demux_004_src8_channel),        //           .channel
		.src8_startofpacket  (cmd_xbar_demux_004_src8_startofpacket),  //           .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_004_src8_endofpacket),    //           .endofpacket
		.src9_ready          (cmd_xbar_demux_004_src9_ready),          //       src9.ready
		.src9_valid          (cmd_xbar_demux_004_src9_valid),          //           .valid
		.src9_data           (cmd_xbar_demux_004_src9_data),           //           .data
		.src9_channel        (cmd_xbar_demux_004_src9_channel),        //           .channel
		.src9_startofpacket  (cmd_xbar_demux_004_src9_startofpacket),  //           .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_004_src9_endofpacket),    //           .endofpacket
		.src10_ready         (cmd_xbar_demux_004_src10_ready),         //      src10.ready
		.src10_valid         (cmd_xbar_demux_004_src10_valid),         //           .valid
		.src10_data          (cmd_xbar_demux_004_src10_data),          //           .data
		.src10_channel       (cmd_xbar_demux_004_src10_channel),       //           .channel
		.src10_startofpacket (cmd_xbar_demux_004_src10_startofpacket), //           .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_004_src10_endofpacket)    //           .endofpacket
	);

	DE0Qsys_rsp_xbar_demux_005 rsp_xbar_demux_005 (
		.clk                (syspll_c0_clk),                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	DE0Qsys_rsp_xbar_demux_005 rsp_xbar_demux_006 (
		.clk                (syspll_c0_clk),                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	DE0Qsys_rsp_xbar_demux_005 rsp_xbar_demux_007 (
		.clk                (syspll_c0_clk),                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	DE0Qsys_rsp_xbar_demux_005 rsp_xbar_demux_008 (
		.clk                (syspll_c0_clk),                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	DE0Qsys_rsp_xbar_demux_005 rsp_xbar_demux_009 (
		.clk                (syspll_c0_clk),                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket)    //          .endofpacket
	);

	DE0Qsys_rsp_xbar_demux_005 rsp_xbar_demux_010 (
		.clk                (syspll_c0_clk),                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_010_src_ready),               //      sink.ready
		.sink_channel       (id_router_010_src_channel),             //          .channel
		.sink_data          (id_router_010_src_data),                //          .data
		.sink_startofpacket (id_router_010_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_010_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_010_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket)    //          .endofpacket
	);

	DE0Qsys_rsp_xbar_demux_005 rsp_xbar_demux_011 (
		.clk                (syspll_c0_clk),                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_011_src_ready),               //      sink.ready
		.sink_channel       (id_router_011_src_channel),             //          .channel
		.sink_data          (id_router_011_src_data),                //          .data
		.sink_startofpacket (id_router_011_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_011_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_011_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_011_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	DE0Qsys_rsp_xbar_demux_005 rsp_xbar_demux_012 (
		.clk                (syspll_c0_clk),                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_012_src_ready),               //      sink.ready
		.sink_channel       (id_router_012_src_channel),             //          .channel
		.sink_data          (id_router_012_src_data),                //          .data
		.sink_startofpacket (id_router_012_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_012_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_012_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_012_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_012_src0_endofpacket)    //          .endofpacket
	);

	DE0Qsys_rsp_xbar_demux_005 rsp_xbar_demux_013 (
		.clk                (syspll_c0_clk),                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_013_src_ready),               //      sink.ready
		.sink_channel       (id_router_013_src_channel),             //          .channel
		.sink_data          (id_router_013_src_data),                //          .data
		.sink_startofpacket (id_router_013_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_013_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_013_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_013_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_013_src0_endofpacket)    //          .endofpacket
	);

	DE0Qsys_rsp_xbar_demux_005 rsp_xbar_demux_014 (
		.clk                (syspll_c0_clk),                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_014_src_ready),               //      sink.ready
		.sink_channel       (id_router_014_src_channel),             //          .channel
		.sink_data          (id_router_014_src_data),                //          .data
		.sink_startofpacket (id_router_014_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_014_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_014_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_014_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_014_src0_endofpacket)    //          .endofpacket
	);

	DE0Qsys_rsp_xbar_demux_005 rsp_xbar_demux_015 (
		.clk                (syspll_c0_clk),                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_015_src_ready),               //      sink.ready
		.sink_channel       (id_router_015_src_channel),             //          .channel
		.sink_data          (id_router_015_src_data),                //          .data
		.sink_startofpacket (id_router_015_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_015_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_015_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_015_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_015_src0_endofpacket)    //          .endofpacket
	);

	DE0Qsys_rsp_xbar_mux_004 rsp_xbar_mux_004 (
		.clk                  (syspll_c0_clk),                         //       clk.clk
		.reset                (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready            (rsp_xbar_mux_004_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_004_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_004_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_004_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_004_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_004_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_005_src0_ready),         //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink0_channel        (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink0_data           (rsp_xbar_demux_005_src0_data),          //          .data
		.sink0_startofpacket  (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_006_src0_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_006_src0_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_007_src0_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_007_src0_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_008_src0_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_008_src0_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_009_src0_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_009_src0_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_009_src0_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_009_src0_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_010_src0_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_010_src0_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_010_src0_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_010_src0_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_011_src0_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_011_src0_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_011_src0_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_011_src0_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_011_src0_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_012_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_012_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_012_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_012_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_012_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_013_src0_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_013_src0_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_013_src0_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_013_src0_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_013_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_014_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_014_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_014_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_014_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_014_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_015_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_015_src0_endofpacket)    //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (61),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (77),
		.IN_PKT_BYTE_CNT_L             (68),
		.IN_PKT_TRANS_COMPRESSED_READ  (62),
		.IN_PKT_BURSTWRAP_H            (80),
		.IN_PKT_BURSTWRAP_L            (78),
		.IN_PKT_BURST_SIZE_H           (83),
		.IN_PKT_BURST_SIZE_L           (81),
		.IN_PKT_RESPONSE_STATUS_H      (105),
		.IN_PKT_RESPONSE_STATUS_L      (104),
		.IN_PKT_TRANS_EXCLUSIVE        (67),
		.IN_PKT_BURST_TYPE_H           (85),
		.IN_PKT_BURST_TYPE_L           (84),
		.IN_ST_DATA_W                  (106),
		.OUT_PKT_ADDR_H                (43),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (59),
		.OUT_PKT_BYTE_CNT_L            (50),
		.OUT_PKT_TRANS_COMPRESSED_READ (44),
		.OUT_PKT_BURST_SIZE_H          (65),
		.OUT_PKT_BURST_SIZE_L          (63),
		.OUT_PKT_RESPONSE_STATUS_H     (87),
		.OUT_PKT_RESPONSE_STATUS_L     (86),
		.OUT_PKT_TRANS_EXCLUSIVE       (49),
		.OUT_PKT_BURST_TYPE_H          (67),
		.OUT_PKT_BURST_TYPE_L          (66),
		.OUT_ST_DATA_W                 (88),
		.ST_CHANNEL_W                  (5),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter (
		.clk                  (syspll_c0_clk),                      //       clk.clk
		.reset                (rst_controller_001_reset_out_reset), // clk_reset.reset
		.in_valid             (cmd_xbar_mux_001_src_valid),         //      sink.valid
		.in_channel           (cmd_xbar_mux_001_src_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_mux_001_src_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_mux_001_src_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_mux_001_src_ready),         //          .ready
		.in_data              (cmd_xbar_mux_001_src_data),          //          .data
		.out_endofpacket      (width_adapter_src_endofpacket),      //       src.endofpacket
		.out_data             (width_adapter_src_data),             //          .data
		.out_channel          (width_adapter_src_channel),          //          .channel
		.out_valid            (width_adapter_src_valid),            //          .valid
		.out_ready            (width_adapter_src_ready),            //          .ready
		.out_startofpacket    (width_adapter_src_startofpacket),    //          .startofpacket
		.in_command_size_data (3'b000)                              // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (43),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (59),
		.IN_PKT_BYTE_CNT_L             (50),
		.IN_PKT_TRANS_COMPRESSED_READ  (44),
		.IN_PKT_BURSTWRAP_H            (62),
		.IN_PKT_BURSTWRAP_L            (60),
		.IN_PKT_BURST_SIZE_H           (65),
		.IN_PKT_BURST_SIZE_L           (63),
		.IN_PKT_RESPONSE_STATUS_H      (87),
		.IN_PKT_RESPONSE_STATUS_L      (86),
		.IN_PKT_TRANS_EXCLUSIVE        (49),
		.IN_PKT_BURST_TYPE_H           (67),
		.IN_PKT_BURST_TYPE_L           (66),
		.IN_ST_DATA_W                  (88),
		.OUT_PKT_ADDR_H                (61),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (77),
		.OUT_PKT_BYTE_CNT_L            (68),
		.OUT_PKT_TRANS_COMPRESSED_READ (62),
		.OUT_PKT_BURST_SIZE_H          (83),
		.OUT_PKT_BURST_SIZE_L          (81),
		.OUT_PKT_RESPONSE_STATUS_H     (105),
		.OUT_PKT_RESPONSE_STATUS_L     (104),
		.OUT_PKT_TRANS_EXCLUSIVE       (67),
		.OUT_PKT_BURST_TYPE_H          (85),
		.OUT_PKT_BURST_TYPE_L          (84),
		.OUT_ST_DATA_W                 (106),
		.ST_CHANNEL_W                  (5),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (1)
	) width_adapter_001 (
		.clk                  (syspll_c0_clk),                       //       clk.clk
		.reset                (rst_controller_001_reset_out_reset),  // clk_reset.reset
		.in_valid             (id_router_001_src_valid),             //      sink.valid
		.in_channel           (id_router_001_src_channel),           //          .channel
		.in_startofpacket     (id_router_001_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_001_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_001_src_ready),             //          .ready
		.in_data              (id_router_001_src_data),              //          .data
		.out_endofpacket      (width_adapter_001_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_001_src_data),          //          .data
		.out_channel          (width_adapter_001_src_channel),       //          .channel
		.out_valid            (width_adapter_001_src_valid),         //          .valid
		.out_ready            (width_adapter_001_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_001_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (106),
		.BITS_PER_SYMBOL     (106),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (5),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser (
		.in_clk            (syspll_c0_clk),                         //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (clk_50m_clk),                           //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_002_src4_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_002_src4_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_002_src4_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_002_src4_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_002_src4_channel),       //              .channel
		.in_data           (cmd_xbar_demux_002_src4_data),          //              .data
		.out_ready         (crosser_out_ready),                     //           out.ready
		.out_valid         (crosser_out_valid),                     //              .valid
		.out_startofpacket (crosser_out_startofpacket),             //              .startofpacket
		.out_endofpacket   (crosser_out_endofpacket),               //              .endofpacket
		.out_channel       (crosser_out_channel),                   //              .channel
		.out_data          (crosser_out_data),                      //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (106),
		.BITS_PER_SYMBOL     (106),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (5),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_001 (
		.in_clk            (clk_50m_clk),                           //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (syspll_c0_clk),                         //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_004_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_004_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_004_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_004_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_004_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_004_src0_data),          //              .data
		.out_ready         (crosser_001_out_ready),                 //           out.ready
		.out_valid         (crosser_001_out_valid),                 //              .valid
		.out_startofpacket (crosser_001_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_001_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_001_out_channel),               //              .channel
		.out_data          (crosser_001_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	DE0Qsys_irq_mapper irq_mapper (
		.clk           (syspll_c0_clk),                      //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.sender_irq    (nios2cpu_d_irq_irq)                  //    sender.irq
	);

endmodule
